

module read_d12 
#(parameter NUM_BITS=10, DEPTH=8)
(

input logic clk,
input logic reset,
input logic [15:10] channel,
input logic [9:0] data,
output logic [15:10] channel_op,
output logic [9:0] data_op,

input logic [7:0] reg1,
input logic [7:0] reg2,
input logic [15:0] concat_data1,

input rst_n,
        //input clk1,
        input rd_en1,
        input wr_en1,
        input [(NUM_BITS-1):0] fifo_in,
        output reg [(NUM_BITS-1):0] fifo_out,
		  input logic [(NUM_BITS+6):0] prevfifo_in, //average
		  input logic [(NUM_BITS+6):0] sum,
		  input logic [(NUM_BITS+6):0] thres,
		  input logic [(NUM_BITS-1):0] Threshold,
        output empty,
        output full,
        output reg [(clogb2(DEPTH)):0] fifo_counter // Able to count more than depth

);


typedef enum logic [63:0] {ch0, ch1, ch2, ch3, ch4 ,ch5, ch6, ch7, ch8, ch9, ch10, ch11, ch12, ch13, ch14, ch15, ch16, ch17, ch18, ch19, ch20, ch21, ch22, ch23, ch24, ch25, ch26, ch27, ch28, ch29, ch30, ch31, ch32, ch33, ch34, ch35, ch36, ch37, ch38, ch39, ch40, ch41, ch42, ch43, ch44, ch45, ch46, ch47, ch48, ch49, ch50, ch51, ch52, ch53, ch54, ch55, ch56,ch57, ch58, ch59, ch60, ch61, ch62, ch63} State;
State currentState, nextState;

always_ff @(posedge clk)
if (reset)
currentState<=ch0;
else currentState<=nextState;

always_comb

case(currentState)

ch0: 
if (channel == 6'b000000) nextState=ch0;
else if (channel ==6'b000001) nextState=ch1;
else if (channel ==6'b000010) nextState=ch2;
else if (channel ==6'b000011) nextState=ch3;
else if (channel ==6'b000100) nextState=ch4;
else if (channel ==6'b000101) nextState=ch5;
else if (channel ==6'b000110) nextState=ch6;
else if (channel ==6'b000111) nextState=ch7;
else if (channel ==6'b001000) nextState=ch8;
else if (channel ==6'b001001) nextState=ch9;
else if (channel ==6'b001010) nextState=ch10;
else if (channel ==6'b001011) nextState=ch11;
else if (channel ==6'b001100) nextState=ch12;
else if (channel ==6'b001101) nextState=ch13;
else if (channel ==6'b001110) nextState=ch14;
else if (channel ==6'b001111) nextState=ch15;
else if (channel ==6'b010000) nextState=ch16;
else if (channel ==6'b010001) nextState=ch17;
else if (channel ==6'b010010) nextState=ch18;
else if (channel ==6'b010011) nextState=ch19;
else if (channel ==6'b010100) nextState=ch20;
else if (channel ==6'b010101) nextState=ch21;
else if (channel ==6'b010110) nextState=ch22;
else if (channel ==6'b010111) nextState=ch23;
else if (channel ==6'b011000) nextState=ch24;
else if (channel ==6'b011001) nextState=ch25;
else if (channel ==6'b011010) nextState=ch26;
else if (channel ==6'b011011) nextState=ch27;
else if (channel ==6'b011100) nextState=ch28;
else if (channel ==6'b011101) nextState=ch29;
else if (channel ==6'b011110) nextState=ch30;
else if (channel ==6'b011111) nextState=ch31;
else if (channel ==6'b100000) nextState=ch32;
else if (channel ==6'b100001) nextState=ch33;
else if (channel ==6'b100010) nextState=ch34;
else if (channel ==6'b100011) nextState=ch35;
else if (channel ==6'b100100) nextState=ch36;
else if (channel ==6'b100101) nextState=ch37;
else if (channel ==6'b100110) nextState=ch38;
else if (channel ==6'b100111) nextState=ch39;
else if (channel ==6'b101000) nextState=ch40;
else if (channel ==6'b101001) nextState=ch41;
else if (channel ==6'b101010) nextState=ch42;
else if (channel ==6'b101011) nextState=ch43;
else if (channel ==6'b101100) nextState=ch44;
else if (channel ==6'b101101) nextState=ch45;
else if (channel ==6'b101110) nextState=ch46;
else if (channel ==6'b101111) nextState=ch47;
else if (channel ==6'b110000) nextState=ch48;
else if (channel ==6'b110001) nextState=ch49;
else if (channel ==6'b110010) nextState=ch50;
else if (channel ==6'b110011) nextState=ch51;
else if (channel ==6'b110100) nextState=ch52;
else if (channel ==6'b110101) nextState=ch53;
else if (channel ==6'b110110) nextState=ch54;
else if (channel ==6'b110111) nextState=ch55;
else if (channel ==6'b111000) nextState=ch56;
else if (channel ==6'b111001) nextState=ch57;
else if (channel ==6'b111010) nextState=ch58;
else if (channel ==6'b111011) nextState=ch59;
else if (channel ==6'b111100) nextState=ch60;
else if (channel ==6'b111101) nextState=ch61;
else if (channel ==6'b111110) nextState=ch62;
else nextState=ch63;


ch1:if (channel ==6'b000001) nextState=ch1;
else if (channel ==6'b000000) nextState=ch0;
else if (channel ==6'b000010) nextState=ch2;
else if (channel ==6'b000011) nextState=ch3;
else if (channel ==6'b000100) nextState=ch4;
else if (channel ==6'b000101) nextState=ch5;
else if (channel ==6'b000110) nextState=ch6;
else if (channel ==6'b000111) nextState=ch7;
else if (channel ==6'b001000) nextState=ch8;
else if (channel ==6'b001001) nextState=ch9;
else if (channel ==6'b001010) nextState=ch10;
else if (channel ==6'b001011) nextState=ch11;
else if (channel ==6'b001100) nextState=ch12;
else if (channel ==6'b001101) nextState=ch13;
else if (channel ==6'b001110) nextState=ch14;
else if (channel ==6'b001111) nextState=ch15;
else if (channel ==6'b010000) nextState=ch16;
else if (channel ==6'b010001) nextState=ch17;
else if (channel ==6'b010010) nextState=ch18;
else if (channel ==6'b010011) nextState=ch19;
else if (channel ==6'b010100) nextState=ch20;
else if (channel ==6'b010101) nextState=ch21;
else if (channel ==6'b010110) nextState=ch22;
else if (channel ==6'b010111) nextState=ch23;
else if (channel ==6'b011000) nextState=ch24;
else if (channel ==6'b011001) nextState=ch25;
else if (channel ==6'b011010) nextState=ch26;
else if (channel ==6'b011011) nextState=ch27;
else if (channel ==6'b011100) nextState=ch28;
else if (channel ==6'b011101) nextState=ch29;
else if (channel ==6'b011110) nextState=ch30;
else if (channel ==6'b011111) nextState=ch31;
else if (channel ==6'b100000) nextState=ch32;
else if (channel ==6'b100001) nextState=ch33;
else if (channel ==6'b100010) nextState=ch34;
else if (channel ==6'b100011) nextState=ch35;
else if (channel ==6'b100100) nextState=ch36;
else if (channel ==6'b100101) nextState=ch37;
else if (channel ==6'b100110) nextState=ch38;
else if (channel ==6'b100111) nextState=ch39;
else if (channel ==6'b101000) nextState=ch40;
else if (channel ==6'b101001) nextState=ch41;
else if (channel ==6'b101010) nextState=ch42;
else if (channel ==6'b101011) nextState=ch43;
else if (channel ==6'b101100) nextState=ch44;
else if (channel ==6'b101101) nextState=ch45;
else if (channel ==6'b101110) nextState=ch46;
else if (channel ==6'b101111) nextState=ch47;
else if (channel ==6'b110000) nextState=ch48;
else if (channel ==6'b110001) nextState=ch49;
else if (channel ==6'b110010) nextState=ch50;
else if (channel ==6'b110011) nextState=ch51;
else if (channel ==6'b110100) nextState=ch52;
else if (channel ==6'b110101) nextState=ch53;
else if (channel ==6'b110110) nextState=ch54;
else if (channel ==6'b110111) nextState=ch55;
else if (channel ==6'b111000) nextState=ch56;
else if (channel ==6'b111001) nextState=ch57;
else if (channel ==6'b111010) nextState=ch58;
else if (channel ==6'b111011) nextState=ch59;
else if (channel ==6'b111100) nextState=ch60;
else if (channel ==6'b111101) nextState=ch61;
else if (channel ==6'b111110) nextState=ch62;
else nextState=ch63;


ch2:if (channel ==6'b000010) nextState=ch2;
else if (channel ==6'b000001) nextState=ch1;
else if (channel ==6'b000000) nextState=ch0;
else if (channel ==6'b000011) nextState=ch3;
else if (channel ==6'b000100) nextState=ch4;
else if (channel ==6'b000101) nextState=ch5;
else if (channel ==6'b000110) nextState=ch6;
else if (channel ==6'b000111) nextState=ch7;
else if (channel ==6'b001000) nextState=ch8;
else if (channel ==6'b001001) nextState=ch9;
else if (channel ==6'b001010) nextState=ch10;
else if (channel ==6'b001011) nextState=ch11;
else if (channel ==6'b001100) nextState=ch12;
else if (channel ==6'b001101) nextState=ch13;
else if (channel ==6'b001110) nextState=ch14;
else if (channel ==6'b001111) nextState=ch15;
else if (channel ==6'b010000) nextState=ch16;
else if (channel ==6'b010001) nextState=ch17;
else if (channel ==6'b010010) nextState=ch18;
else if (channel ==6'b010011) nextState=ch19;
else if (channel ==6'b010100) nextState=ch20;
else if (channel ==6'b010101) nextState=ch21;
else if (channel ==6'b010110) nextState=ch22;
else if (channel ==6'b010111) nextState=ch23;
else if (channel ==6'b011000) nextState=ch24;
else if (channel ==6'b011001) nextState=ch25;
else if (channel ==6'b011010) nextState=ch26;
else if (channel ==6'b011011) nextState=ch27;
else if (channel ==6'b011100) nextState=ch28;
else if (channel ==6'b011101) nextState=ch29;
else if (channel ==6'b011110) nextState=ch30;
else if (channel ==6'b011111) nextState=ch31;
else if (channel ==6'b100000) nextState=ch32;
else if (channel ==6'b100001) nextState=ch33;
else if (channel ==6'b100010) nextState=ch34;
else if (channel ==6'b100011) nextState=ch35;
else if (channel ==6'b100100) nextState=ch36;
else if (channel ==6'b100101) nextState=ch37;
else if (channel ==6'b100110) nextState=ch38;
else if (channel ==6'b100111) nextState=ch39;
else if (channel ==6'b101000) nextState=ch40;
else if (channel ==6'b101001) nextState=ch41;
else if (channel ==6'b101010) nextState=ch42;
else if (channel ==6'b101011) nextState=ch43;
else if (channel ==6'b101100) nextState=ch44;
else if (channel ==6'b101101) nextState=ch45;
else if (channel ==6'b101110) nextState=ch46;
else if (channel ==6'b101111) nextState=ch47;
else if (channel ==6'b110000) nextState=ch48;
else if (channel ==6'b110001) nextState=ch49;
else if (channel ==6'b110010) nextState=ch50;
else if (channel ==6'b110011) nextState=ch51;
else if (channel ==6'b110100) nextState=ch52;
else if (channel ==6'b110101) nextState=ch53;
else if (channel ==6'b110110) nextState=ch54;
else if (channel ==6'b110111) nextState=ch55;
else if (channel ==6'b111000) nextState=ch56;
else if (channel ==6'b111001) nextState=ch57;
else if (channel ==6'b111010) nextState=ch58;
else if (channel ==6'b111011) nextState=ch59;
else if (channel ==6'b111100) nextState=ch60;
else if (channel ==6'b111101) nextState=ch61;
else if (channel ==6'b111110) nextState=ch62;
else nextState=ch63;

ch3:if (channel ==6'b000011) nextState=ch3;
else if (channel ==6'b000001) nextState=ch1;
else if (channel ==6'b000010) nextState=ch2;
else if (channel ==6'b000000) nextState=ch0;
else if (channel ==6'b000100) nextState=ch4;
else if (channel ==6'b000101) nextState=ch5;
else if (channel ==6'b000110) nextState=ch6;
else if (channel ==6'b000111) nextState=ch7;
else if (channel ==6'b001000) nextState=ch8;
else if (channel ==6'b001001) nextState=ch9;
else if (channel ==6'b001010) nextState=ch10;
else if (channel ==6'b001011) nextState=ch11;
else if (channel ==6'b001100) nextState=ch12;
else if (channel ==6'b001101) nextState=ch13;
else if (channel ==6'b001110) nextState=ch14;
else if (channel ==6'b001111) nextState=ch15;
else if (channel ==6'b010000) nextState=ch16;
else if (channel ==6'b010001) nextState=ch17;
else if (channel ==6'b010010) nextState=ch18;
else if (channel ==6'b010011) nextState=ch19;
else if (channel ==6'b010100) nextState=ch20;
else if (channel ==6'b010101) nextState=ch21;
else if (channel ==6'b010110) nextState=ch22;
else if (channel ==6'b010111) nextState=ch23;
else if (channel ==6'b011000) nextState=ch24;
else if (channel ==6'b011001) nextState=ch25;
else if (channel ==6'b011010) nextState=ch26;
else if (channel ==6'b011011) nextState=ch27;
else if (channel ==6'b011100) nextState=ch28;
else if (channel ==6'b011101) nextState=ch29;
else if (channel ==6'b011110) nextState=ch30;
else if (channel ==6'b011111) nextState=ch31;
else if (channel ==6'b100000) nextState=ch32;
else if (channel ==6'b100001) nextState=ch33;
else if (channel ==6'b100010) nextState=ch34;
else if (channel ==6'b100011) nextState=ch35;
else if (channel ==6'b100100) nextState=ch36;
else if (channel ==6'b100101) nextState=ch37;
else if (channel ==6'b100110) nextState=ch38;
else if (channel ==6'b100111) nextState=ch39;
else if (channel ==6'b101000) nextState=ch40;
else if (channel ==6'b101001) nextState=ch41;
else if (channel ==6'b101010) nextState=ch42;
else if (channel ==6'b101011) nextState=ch43;
else if (channel ==6'b101100) nextState=ch44;
else if (channel ==6'b101101) nextState=ch45;
else if (channel ==6'b101110) nextState=ch46;
else if (channel ==6'b101111) nextState=ch47;
else if (channel ==6'b110000) nextState=ch48;
else if (channel ==6'b110001) nextState=ch49;
else if (channel ==6'b110010) nextState=ch50;
else if (channel ==6'b110011) nextState=ch51;
else if (channel ==6'b110100) nextState=ch52;
else if (channel ==6'b110101) nextState=ch53;
else if (channel ==6'b110110) nextState=ch54;
else if (channel ==6'b110111) nextState=ch55;
else if (channel ==6'b111000) nextState=ch56;
else if (channel ==6'b111001) nextState=ch57;
else if (channel ==6'b111010) nextState=ch58;
else if (channel ==6'b111011) nextState=ch59;
else if (channel ==6'b111100) nextState=ch60;
else if (channel ==6'b111101) nextState=ch61;
else if (channel ==6'b111110) nextState=ch62;
else nextState=ch63;



ch4:if (channel ==6'b000100) nextState=ch4;
else if (channel ==6'b000001) nextState=ch1;
else if (channel ==6'b000010) nextState=ch2;
else if (channel ==6'b000011) nextState=ch3;
else if (channel ==6'b000000) nextState=ch0;
else if (channel ==6'b000101) nextState=ch5;
else if (channel ==6'b000110) nextState=ch6;
else if (channel ==6'b000111) nextState=ch7;
else if (channel ==6'b001000) nextState=ch8;
else if (channel ==6'b001001) nextState=ch9;
else if (channel ==6'b001010) nextState=ch10;
else if (channel ==6'b001011) nextState=ch11;
else if (channel ==6'b001100) nextState=ch12;
else if (channel ==6'b001101) nextState=ch13;
else if (channel ==6'b001110) nextState=ch14;
else if (channel ==6'b001111) nextState=ch15;
else if (channel ==6'b010000) nextState=ch16;
else if (channel ==6'b010001) nextState=ch17;
else if (channel ==6'b010010) nextState=ch18;
else if (channel ==6'b010011) nextState=ch19;
else if (channel ==6'b010100) nextState=ch20;
else if (channel ==6'b010101) nextState=ch21;
else if (channel ==6'b010110) nextState=ch22;
else if (channel ==6'b010111) nextState=ch23;
else if (channel ==6'b011000) nextState=ch24;
else if (channel ==6'b011001) nextState=ch25;
else if (channel ==6'b011010) nextState=ch26;
else if (channel ==6'b011011) nextState=ch27;
else if (channel ==6'b011100) nextState=ch28;
else if (channel ==6'b011101) nextState=ch29;
else if (channel ==6'b011110) nextState=ch30;
else if (channel ==6'b011111) nextState=ch31;
else if (channel ==6'b100000) nextState=ch32;
else if (channel ==6'b100001) nextState=ch33;
else if (channel ==6'b100010) nextState=ch34;
else if (channel ==6'b100011) nextState=ch35;
else if (channel ==6'b100100) nextState=ch36;
else if (channel ==6'b100101) nextState=ch37;
else if (channel ==6'b100110) nextState=ch38;
else if (channel ==6'b100111) nextState=ch39;
else if (channel ==6'b101000) nextState=ch40;
else if (channel ==6'b101001) nextState=ch41;
else if (channel ==6'b101010) nextState=ch42;
else if (channel ==6'b101011) nextState=ch43;
else if (channel ==6'b101100) nextState=ch44;
else if (channel ==6'b101101) nextState=ch45;
else if (channel ==6'b101110) nextState=ch46;
else if (channel ==6'b101111) nextState=ch47;
else if (channel ==6'b110000) nextState=ch48;
else if (channel ==6'b110001) nextState=ch49;
else if (channel ==6'b110010) nextState=ch50;
else if (channel ==6'b110011) nextState=ch51;
else if (channel ==6'b110100) nextState=ch52;
else if (channel ==6'b110101) nextState=ch53;
else if (channel ==6'b110110) nextState=ch54;
else if (channel ==6'b110111) nextState=ch55;
else if (channel ==6'b111000) nextState=ch56;
else if (channel ==6'b111001) nextState=ch57;
else if (channel ==6'b111010) nextState=ch58;
else if (channel ==6'b111011) nextState=ch59;
else if (channel ==6'b111100) nextState=ch60;
else if (channel ==6'b111101) nextState=ch61;
else if (channel ==6'b111110) nextState=ch62;
else nextState=ch63;



ch5:if (channel ==6'b000101) nextState=ch5;
else if (channel ==6'b000001) nextState=ch1;
else if (channel ==6'b000010) nextState=ch2;
else if (channel ==6'b000011) nextState=ch3;
else if (channel ==6'b000100) nextState=ch4;
else if (channel ==6'b000000) nextState=ch0;
else if (channel ==6'b000110) nextState=ch6;
else if (channel ==6'b000111) nextState=ch7;
else if (channel ==6'b001000) nextState=ch8;
else if (channel ==6'b001001) nextState=ch9;
else if (channel ==6'b001010) nextState=ch10;
else if (channel ==6'b001011) nextState=ch11;
else if (channel ==6'b001100) nextState=ch12;
else if (channel ==6'b001101) nextState=ch13;
else if (channel ==6'b001110) nextState=ch14;
else if (channel ==6'b001111) nextState=ch15;
else if (channel ==6'b010000) nextState=ch16;
else if (channel ==6'b010001) nextState=ch17;
else if (channel ==6'b010010) nextState=ch18;
else if (channel ==6'b010011) nextState=ch19;
else if (channel ==6'b010100) nextState=ch20;
else if (channel ==6'b010101) nextState=ch21;
else if (channel ==6'b010110) nextState=ch22;
else if (channel ==6'b010111) nextState=ch23;
else if (channel ==6'b011000) nextState=ch24;
else if (channel ==6'b011001) nextState=ch25;
else if (channel ==6'b011010) nextState=ch26;
else if (channel ==6'b011011) nextState=ch27;
else if (channel ==6'b011100) nextState=ch28;
else if (channel ==6'b011101) nextState=ch29;
else if (channel ==6'b011110) nextState=ch30;
else if (channel ==6'b011111) nextState=ch31;
else if (channel ==6'b100000) nextState=ch32;
else if (channel ==6'b100001) nextState=ch33;
else if (channel ==6'b100010) nextState=ch34;
else if (channel ==6'b100011) nextState=ch35;
else if (channel ==6'b100100) nextState=ch36;
else if (channel ==6'b100101) nextState=ch37;
else if (channel ==6'b100110) nextState=ch38;
else if (channel ==6'b100111) nextState=ch39;
else if (channel ==6'b101000) nextState=ch40;
else if (channel ==6'b101001) nextState=ch41;
else if (channel ==6'b101010) nextState=ch42;
else if (channel ==6'b101011) nextState=ch43;
else if (channel ==6'b101100) nextState=ch44;
else if (channel ==6'b101101) nextState=ch45;
else if (channel ==6'b101110) nextState=ch46;
else if (channel ==6'b101111) nextState=ch47;
else if (channel ==6'b110000) nextState=ch48;
else if (channel ==6'b110001) nextState=ch49;
else if (channel ==6'b110010) nextState=ch50;
else if (channel ==6'b110011) nextState=ch51;
else if (channel ==6'b110100) nextState=ch52;
else if (channel ==6'b110101) nextState=ch53;
else if (channel ==6'b110110) nextState=ch54;
else if (channel ==6'b110111) nextState=ch55;
else if (channel ==6'b111000) nextState=ch56;
else if (channel ==6'b111001) nextState=ch57;
else if (channel ==6'b111010) nextState=ch58;
else if (channel ==6'b111011) nextState=ch59;
else if (channel ==6'b111100) nextState=ch60;
else if (channel ==6'b111101) nextState=ch61;
else if (channel ==6'b111110) nextState=ch62;
else nextState=ch63;



ch6:if (channel ==6'b000110) nextState=ch6;
else if (channel ==6'b000001) nextState=ch1;
else if (channel ==6'b000010) nextState=ch2;
else if (channel ==6'b000011) nextState=ch3;
else if (channel ==6'b000100) nextState=ch4;
else if (channel ==6'b000101) nextState=ch5;
else if (channel ==6'b000000) nextState=ch0;
else if (channel ==6'b000111) nextState=ch7;
else if (channel ==6'b001000) nextState=ch8;
else if (channel ==6'b001001) nextState=ch9;
else if (channel ==6'b001010) nextState=ch10;
else if (channel ==6'b001011) nextState=ch11;
else if (channel ==6'b001100) nextState=ch12;
else if (channel ==6'b001101) nextState=ch13;
else if (channel ==6'b001110) nextState=ch14;
else if (channel ==6'b001111) nextState=ch15;
else if (channel ==6'b010000) nextState=ch16;
else if (channel ==6'b010001) nextState=ch17;
else if (channel ==6'b010010) nextState=ch18;
else if (channel ==6'b010011) nextState=ch19;
else if (channel ==6'b010100) nextState=ch20;
else if (channel ==6'b010101) nextState=ch21;
else if (channel ==6'b010110) nextState=ch22;
else if (channel ==6'b010111) nextState=ch23;
else if (channel ==6'b011000) nextState=ch24;
else if (channel ==6'b011001) nextState=ch25;
else if (channel ==6'b011010) nextState=ch26;
else if (channel ==6'b011011) nextState=ch27;
else if (channel ==6'b011100) nextState=ch28;
else if (channel ==6'b011101) nextState=ch29;
else if (channel ==6'b011110) nextState=ch30;
else if (channel ==6'b011111) nextState=ch31;
else if (channel ==6'b100000) nextState=ch32;
else if (channel ==6'b100001) nextState=ch33;
else if (channel ==6'b100010) nextState=ch34;
else if (channel ==6'b100011) nextState=ch35;
else if (channel ==6'b100100) nextState=ch36;
else if (channel ==6'b100101) nextState=ch37;
else if (channel ==6'b100110) nextState=ch38;
else if (channel ==6'b100111) nextState=ch39;
else if (channel ==6'b101000) nextState=ch40;
else if (channel ==6'b101001) nextState=ch41;
else if (channel ==6'b101010) nextState=ch42;
else if (channel ==6'b101011) nextState=ch43;
else if (channel ==6'b101100) nextState=ch44;
else if (channel ==6'b101101) nextState=ch45;
else if (channel ==6'b101110) nextState=ch46;
else if (channel ==6'b101111) nextState=ch47;
else if (channel ==6'b110000) nextState=ch48;
else if (channel ==6'b110001) nextState=ch49;
else if (channel ==6'b110010) nextState=ch50;
else if (channel ==6'b110011) nextState=ch51;
else if (channel ==6'b110100) nextState=ch52;
else if (channel ==6'b110101) nextState=ch53;
else if (channel ==6'b110110) nextState=ch54;
else if (channel ==6'b110111) nextState=ch55;
else if (channel ==6'b111000) nextState=ch56;
else if (channel ==6'b111001) nextState=ch57;
else if (channel ==6'b111010) nextState=ch58;
else if (channel ==6'b111011) nextState=ch59;
else if (channel ==6'b111100) nextState=ch60;
else if (channel ==6'b111101) nextState=ch61;
else if (channel ==6'b111110) nextState=ch62;
else nextState=ch63;



ch7:if (channel ==6'b000111) nextState=ch7;
else if (channel ==6'b000001) nextState=ch1;
else if (channel ==6'b000010) nextState=ch2;
else if (channel ==6'b000011) nextState=ch3;
else if (channel ==6'b000100) nextState=ch4;
else if (channel ==6'b000101) nextState=ch5;
else if (channel ==6'b000110) nextState=ch6;
else if (channel ==6'b000000) nextState=ch0;
else if (channel ==6'b001000) nextState=ch8;
else if (channel ==6'b001001) nextState=ch9;
else if (channel ==6'b001010) nextState=ch10;
else if (channel ==6'b001011) nextState=ch11;
else if (channel ==6'b001100) nextState=ch12;
else if (channel ==6'b001101) nextState=ch13;
else if (channel ==6'b001110) nextState=ch14;
else if (channel ==6'b001111) nextState=ch15;
else if (channel ==6'b010000) nextState=ch16;
else if (channel ==6'b010001) nextState=ch17;
else if (channel ==6'b010010) nextState=ch18;
else if (channel ==6'b010011) nextState=ch19;
else if (channel ==6'b010100) nextState=ch20;
else if (channel ==6'b010101) nextState=ch21;
else if (channel ==6'b010110) nextState=ch22;
else if (channel ==6'b010111) nextState=ch23;
else if (channel ==6'b011000) nextState=ch24;
else if (channel ==6'b011001) nextState=ch25;
else if (channel ==6'b011010) nextState=ch26;
else if (channel ==6'b011011) nextState=ch27;
else if (channel ==6'b011100) nextState=ch28;
else if (channel ==6'b011101) nextState=ch29;
else if (channel ==6'b011110) nextState=ch30;
else if (channel ==6'b011111) nextState=ch31;
else if (channel ==6'b100000) nextState=ch32;
else if (channel ==6'b100001) nextState=ch33;
else if (channel ==6'b100010) nextState=ch34;
else if (channel ==6'b100011) nextState=ch35;
else if (channel ==6'b100100) nextState=ch36;
else if (channel ==6'b100101) nextState=ch37;
else if (channel ==6'b100110) nextState=ch38;
else if (channel ==6'b100111) nextState=ch39;
else if (channel ==6'b101000) nextState=ch40;
else if (channel ==6'b101001) nextState=ch41;
else if (channel ==6'b101010) nextState=ch42;
else if (channel ==6'b101011) nextState=ch43;
else if (channel ==6'b101100) nextState=ch44;
else if (channel ==6'b101101) nextState=ch45;
else if (channel ==6'b101110) nextState=ch46;
else if (channel ==6'b101111) nextState=ch47;
else if (channel ==6'b110000) nextState=ch48;
else if (channel ==6'b110001) nextState=ch49;
else if (channel ==6'b110010) nextState=ch50;
else if (channel ==6'b110011) nextState=ch51;
else if (channel ==6'b110100) nextState=ch52;
else if (channel ==6'b110101) nextState=ch53;
else if (channel ==6'b110110) nextState=ch54;
else if (channel ==6'b110111) nextState=ch55;
else if (channel ==6'b111000) nextState=ch56;
else if (channel ==6'b111001) nextState=ch57;
else if (channel ==6'b111010) nextState=ch58;
else if (channel ==6'b111011) nextState=ch59;
else if (channel ==6'b111100) nextState=ch60;
else if (channel ==6'b111101) nextState=ch61;
else if (channel ==6'b111110) nextState=ch62;
else nextState=ch63;



ch8:if (channel ==6'b001000) nextState=ch8;
else if (channel ==6'b000001) nextState=ch1;
else if (channel ==6'b000010) nextState=ch2;
else if (channel ==6'b000011) nextState=ch3;
else if (channel ==6'b000100) nextState=ch4;
else if (channel ==6'b000101) nextState=ch5;
else if (channel ==6'b000110) nextState=ch6;
else if (channel ==6'b000111) nextState=ch7;
else if (channel ==6'b000000) nextState=ch0;
else if (channel ==6'b001001) nextState=ch9;
else if (channel ==6'b001010) nextState=ch10;
else if (channel ==6'b001011) nextState=ch11;
else if (channel ==6'b001100) nextState=ch12;
else if (channel ==6'b001101) nextState=ch13;
else if (channel ==6'b001110) nextState=ch14;
else if (channel ==6'b001111) nextState=ch15;
else if (channel ==6'b010000) nextState=ch16;
else if (channel ==6'b010001) nextState=ch17;
else if (channel ==6'b010010) nextState=ch18;
else if (channel ==6'b010011) nextState=ch19;
else if (channel ==6'b010100) nextState=ch20;
else if (channel ==6'b010101) nextState=ch21;
else if (channel ==6'b010110) nextState=ch22;
else if (channel ==6'b010111) nextState=ch23;
else if (channel ==6'b011000) nextState=ch24;
else if (channel ==6'b011001) nextState=ch25;
else if (channel ==6'b011010) nextState=ch26;
else if (channel ==6'b011011) nextState=ch27;
else if (channel ==6'b011100) nextState=ch28;
else if (channel ==6'b011101) nextState=ch29;
else if (channel ==6'b011110) nextState=ch30;
else if (channel ==6'b011111) nextState=ch31;
else if (channel ==6'b100000) nextState=ch32;
else if (channel ==6'b100001) nextState=ch33;
else if (channel ==6'b100010) nextState=ch34;
else if (channel ==6'b100011) nextState=ch35;
else if (channel ==6'b100100) nextState=ch36;
else if (channel ==6'b100101) nextState=ch37;
else if (channel ==6'b100110) nextState=ch38;
else if (channel ==6'b100111) nextState=ch39;
else if (channel ==6'b101000) nextState=ch40;
else if (channel ==6'b101001) nextState=ch41;
else if (channel ==6'b101010) nextState=ch42;
else if (channel ==6'b101011) nextState=ch43;
else if (channel ==6'b101100) nextState=ch44;
else if (channel ==6'b101101) nextState=ch45;
else if (channel ==6'b101110) nextState=ch46;
else if (channel ==6'b101111) nextState=ch47;
else if (channel ==6'b110000) nextState=ch48;
else if (channel ==6'b110001) nextState=ch49;
else if (channel ==6'b110010) nextState=ch50;
else if (channel ==6'b110011) nextState=ch51;
else if (channel ==6'b110100) nextState=ch52;
else if (channel ==6'b110101) nextState=ch53;
else if (channel ==6'b110110) nextState=ch54;
else if (channel ==6'b110111) nextState=ch55;
else if (channel ==6'b111000) nextState=ch56;
else if (channel ==6'b111001) nextState=ch57;
else if (channel ==6'b111010) nextState=ch58;
else if (channel ==6'b111011) nextState=ch59;
else if (channel ==6'b111100) nextState=ch60;
else if (channel ==6'b111101) nextState=ch61;
else if (channel ==6'b111110) nextState=ch62;
else nextState=ch63;



ch9:if (channel ==6'b001001) nextState=ch9;
else if (channel ==6'b000001) nextState=ch1;
else if (channel ==6'b000010) nextState=ch2;
else if (channel ==6'b000011) nextState=ch3;
else if (channel ==6'b000100) nextState=ch4;
else if (channel ==6'b000101) nextState=ch5;
else if (channel ==6'b000110) nextState=ch6;
else if (channel ==6'b000111) nextState=ch7;
else if (channel ==6'b001000) nextState=ch8;
else if (channel ==6'b000000) nextState=ch0;
else if (channel ==6'b001010) nextState=ch10;
else if (channel ==6'b001011) nextState=ch11;
else if (channel ==6'b001100) nextState=ch12;
else if (channel ==6'b001101) nextState=ch13;
else if (channel ==6'b001110) nextState=ch14;
else if (channel ==6'b001111) nextState=ch15;
else if (channel ==6'b010000) nextState=ch16;
else if (channel ==6'b010001) nextState=ch17;
else if (channel ==6'b010010) nextState=ch18;
else if (channel ==6'b010011) nextState=ch19;
else if (channel ==6'b010100) nextState=ch20;
else if (channel ==6'b010101) nextState=ch21;
else if (channel ==6'b010110) nextState=ch22;
else if (channel ==6'b010111) nextState=ch23;
else if (channel ==6'b011000) nextState=ch24;
else if (channel ==6'b011001) nextState=ch25;
else if (channel ==6'b011010) nextState=ch26;
else if (channel ==6'b011011) nextState=ch27;
else if (channel ==6'b011100) nextState=ch28;
else if (channel ==6'b011101) nextState=ch29;
else if (channel ==6'b011110) nextState=ch30;
else if (channel ==6'b011111) nextState=ch31;
else if (channel ==6'b100000) nextState=ch32;
else if (channel ==6'b100001) nextState=ch33;
else if (channel ==6'b100010) nextState=ch34;
else if (channel ==6'b100011) nextState=ch35;
else if (channel ==6'b100100) nextState=ch36;
else if (channel ==6'b100101) nextState=ch37;
else if (channel ==6'b100110) nextState=ch38;
else if (channel ==6'b100111) nextState=ch39;
else if (channel ==6'b101000) nextState=ch40;
else if (channel ==6'b101001) nextState=ch41;
else if (channel ==6'b101010) nextState=ch42;
else if (channel ==6'b101011) nextState=ch43;
else if (channel ==6'b101100) nextState=ch44;
else if (channel ==6'b101101) nextState=ch45;
else if (channel ==6'b101110) nextState=ch46;
else if (channel ==6'b101111) nextState=ch47;
else if (channel ==6'b110000) nextState=ch48;
else if (channel ==6'b110001) nextState=ch49;
else if (channel ==6'b110010) nextState=ch50;
else if (channel ==6'b110011) nextState=ch51;
else if (channel ==6'b110100) nextState=ch52;
else if (channel ==6'b110101) nextState=ch53;
else if (channel ==6'b110110) nextState=ch54;
else if (channel ==6'b110111) nextState=ch55;
else if (channel ==6'b111000) nextState=ch56;
else if (channel ==6'b111001) nextState=ch57;
else if (channel ==6'b111010) nextState=ch58;
else if (channel ==6'b111011) nextState=ch59;
else if (channel ==6'b111100) nextState=ch60;
else if (channel ==6'b111101) nextState=ch61;
else if (channel ==6'b111110) nextState=ch62;
else nextState=ch63;


ch10:if (channel ==6'b001010) nextState=ch10;
else if (channel ==6'b000001) nextState=ch1;
else if (channel ==6'b000010) nextState=ch2;
else if (channel ==6'b000011) nextState=ch3;
else if (channel ==6'b000100) nextState=ch4;
else if (channel ==6'b000101) nextState=ch5;
else if (channel ==6'b000110) nextState=ch6;
else if (channel ==6'b000111) nextState=ch7;
else if (channel ==6'b001000) nextState=ch8;
else if (channel ==6'b001001) nextState=ch9;
else if (channel ==6'b000000) nextState=ch0;
else if (channel ==6'b001011) nextState=ch11;
else if (channel ==6'b001100) nextState=ch12;
else if (channel ==6'b001101) nextState=ch13;
else if (channel ==6'b001110) nextState=ch14;
else if (channel ==6'b001111) nextState=ch15;
else if (channel ==6'b010000) nextState=ch16;
else if (channel ==6'b010001) nextState=ch17;
else if (channel ==6'b010010) nextState=ch18;
else if (channel ==6'b010011) nextState=ch19;
else if (channel ==6'b010100) nextState=ch20;
else if (channel ==6'b010101) nextState=ch21;
else if (channel ==6'b010110) nextState=ch22;
else if (channel ==6'b010111) nextState=ch23;
else if (channel ==6'b011000) nextState=ch24;
else if (channel ==6'b011001) nextState=ch25;
else if (channel ==6'b011010) nextState=ch26;
else if (channel ==6'b011011) nextState=ch27;
else if (channel ==6'b011100) nextState=ch28;
else if (channel ==6'b011101) nextState=ch29;
else if (channel ==6'b011110) nextState=ch30;
else if (channel ==6'b011111) nextState=ch31;
else if (channel ==6'b100000) nextState=ch32;
else if (channel ==6'b100001) nextState=ch33;
else if (channel ==6'b100010) nextState=ch34;
else if (channel ==6'b100011) nextState=ch35;
else if (channel ==6'b100100) nextState=ch36;
else if (channel ==6'b100101) nextState=ch37;
else if (channel ==6'b100110) nextState=ch38;
else if (channel ==6'b100111) nextState=ch39;
else if (channel ==6'b101000) nextState=ch40;
else if (channel ==6'b101001) nextState=ch41;
else if (channel ==6'b101010) nextState=ch42;
else if (channel ==6'b101011) nextState=ch43;
else if (channel ==6'b101100) nextState=ch44;
else if (channel ==6'b101101) nextState=ch45;
else if (channel ==6'b101110) nextState=ch46;
else if (channel ==6'b101111) nextState=ch47;
else if (channel ==6'b110000) nextState=ch48;
else if (channel ==6'b110001) nextState=ch49;
else if (channel ==6'b110010) nextState=ch50;
else if (channel ==6'b110011) nextState=ch51;
else if (channel ==6'b110100) nextState=ch52;
else if (channel ==6'b110101) nextState=ch53;
else if (channel ==6'b110110) nextState=ch54;
else if (channel ==6'b110111) nextState=ch55;
else if (channel ==6'b111000) nextState=ch56;
else if (channel ==6'b111001) nextState=ch57;
else if (channel ==6'b111010) nextState=ch58;
else if (channel ==6'b111011) nextState=ch59;
else if (channel ==6'b111100) nextState=ch60;
else if (channel ==6'b111101) nextState=ch61;
else if (channel ==6'b111110) nextState=ch62;
else nextState=ch63;

ch11:if (channel ==6'b001011) nextState=ch11;
else if (channel ==6'b000001) nextState=ch1;
else if (channel ==6'b000010) nextState=ch2;
else if (channel ==6'b000011) nextState=ch3;
else if (channel ==6'b000100) nextState=ch4;
else if (channel ==6'b000101) nextState=ch5;
else if (channel ==6'b000110) nextState=ch6;
else if (channel ==6'b000111) nextState=ch7;
else if (channel ==6'b001000) nextState=ch8;
else if (channel ==6'b001001) nextState=ch9;
else if (channel ==6'b001010) nextState=ch10;
else if (channel ==6'b000000) nextState=ch0;
else if (channel ==6'b001100) nextState=ch12;
else if (channel ==6'b001101) nextState=ch13;
else if (channel ==6'b001110) nextState=ch14;
else if (channel ==6'b001111) nextState=ch15;
else if (channel ==6'b010000) nextState=ch16;
else if (channel ==6'b010001) nextState=ch17;
else if (channel ==6'b010010) nextState=ch18;
else if (channel ==6'b010011) nextState=ch19;
else if (channel ==6'b010100) nextState=ch20;
else if (channel ==6'b010101) nextState=ch21;
else if (channel ==6'b010110) nextState=ch22;
else if (channel ==6'b010111) nextState=ch23;
else if (channel ==6'b011000) nextState=ch24;
else if (channel ==6'b011001) nextState=ch25;
else if (channel ==6'b011010) nextState=ch26;
else if (channel ==6'b011011) nextState=ch27;
else if (channel ==6'b011100) nextState=ch28;
else if (channel ==6'b011101) nextState=ch29;
else if (channel ==6'b011110) nextState=ch30;
else if (channel ==6'b011111) nextState=ch31;
else if (channel ==6'b100000) nextState=ch32;
else if (channel ==6'b100001) nextState=ch33;
else if (channel ==6'b100010) nextState=ch34;
else if (channel ==6'b100011) nextState=ch35;
else if (channel ==6'b100100) nextState=ch36;
else if (channel ==6'b100101) nextState=ch37;
else if (channel ==6'b100110) nextState=ch38;
else if (channel ==6'b100111) nextState=ch39;
else if (channel ==6'b101000) nextState=ch40;
else if (channel ==6'b101001) nextState=ch41;
else if (channel ==6'b101010) nextState=ch42;
else if (channel ==6'b101011) nextState=ch43;
else if (channel ==6'b101100) nextState=ch44;
else if (channel ==6'b101101) nextState=ch45;
else if (channel ==6'b101110) nextState=ch46;
else if (channel ==6'b101111) nextState=ch47;
else if (channel ==6'b110000) nextState=ch48;
else if (channel ==6'b110001) nextState=ch49;
else if (channel ==6'b110010) nextState=ch50;
else if (channel ==6'b110011) nextState=ch51;
else if (channel ==6'b110100) nextState=ch52;
else if (channel ==6'b110101) nextState=ch53;
else if (channel ==6'b110110) nextState=ch54;
else if (channel ==6'b110111) nextState=ch55;
else if (channel ==6'b111000) nextState=ch56;
else if (channel ==6'b111001) nextState=ch57;
else if (channel ==6'b111010) nextState=ch58;
else if (channel ==6'b111011) nextState=ch59;
else if (channel ==6'b111100) nextState=ch60;
else if (channel ==6'b111101) nextState=ch61;
else if (channel ==6'b111110) nextState=ch62;
else nextState=ch63;


ch12:if (channel ==6'b001100) nextState=ch12;
else if (channel ==6'b000001) nextState=ch1;
else if (channel ==6'b000010) nextState=ch2;
else if (channel ==6'b000011) nextState=ch3;
else if (channel ==6'b000100) nextState=ch4;
else if (channel ==6'b000101) nextState=ch5;
else if (channel ==6'b000110) nextState=ch6;
else if (channel ==6'b000111) nextState=ch7;
else if (channel ==6'b001000) nextState=ch8;
else if (channel ==6'b001001) nextState=ch9;
else if (channel ==6'b001010) nextState=ch10;
else if (channel ==6'b001011) nextState=ch11;
else if (channel ==6'b000000) nextState=ch0;
else if (channel ==6'b001101) nextState=ch13;
else if (channel ==6'b001110) nextState=ch14;
else if (channel ==6'b001111) nextState=ch15;
else if (channel ==6'b010000) nextState=ch16;
else if (channel ==6'b010001) nextState=ch17;
else if (channel ==6'b010010) nextState=ch18;
else if (channel ==6'b010011) nextState=ch19;
else if (channel ==6'b010100) nextState=ch20;
else if (channel ==6'b010101) nextState=ch21;
else if (channel ==6'b010110) nextState=ch22;
else if (channel ==6'b010111) nextState=ch23;
else if (channel ==6'b011000) nextState=ch24;
else if (channel ==6'b011001) nextState=ch25;
else if (channel ==6'b011010) nextState=ch26;
else if (channel ==6'b011011) nextState=ch27;
else if (channel ==6'b011100) nextState=ch28;
else if (channel ==6'b011101) nextState=ch29;
else if (channel ==6'b011110) nextState=ch30;
else if (channel ==6'b011111) nextState=ch31;
else if (channel ==6'b100000) nextState=ch32;
else if (channel ==6'b100001) nextState=ch33;
else if (channel ==6'b100010) nextState=ch34;
else if (channel ==6'b100011) nextState=ch35;
else if (channel ==6'b100100) nextState=ch36;
else if (channel ==6'b100101) nextState=ch37;
else if (channel ==6'b100110) nextState=ch38;
else if (channel ==6'b100111) nextState=ch39;
else if (channel ==6'b101000) nextState=ch40;
else if (channel ==6'b101001) nextState=ch41;
else if (channel ==6'b101010) nextState=ch42;
else if (channel ==6'b101011) nextState=ch43;
else if (channel ==6'b101100) nextState=ch44;
else if (channel ==6'b101101) nextState=ch45;
else if (channel ==6'b101110) nextState=ch46;
else if (channel ==6'b101111) nextState=ch47;
else if (channel ==6'b110000) nextState=ch48;
else if (channel ==6'b110001) nextState=ch49;
else if (channel ==6'b110010) nextState=ch50;
else if (channel ==6'b110011) nextState=ch51;
else if (channel ==6'b110100) nextState=ch52;
else if (channel ==6'b110101) nextState=ch53;
else if (channel ==6'b110110) nextState=ch54;
else if (channel ==6'b110111) nextState=ch55;
else if (channel ==6'b111000) nextState=ch56;
else if (channel ==6'b111001) nextState=ch57;
else if (channel ==6'b111010) nextState=ch58;
else if (channel ==6'b111011) nextState=ch59;
else if (channel ==6'b111100) nextState=ch60;
else if (channel ==6'b111101) nextState=ch61;
else if (channel ==6'b111110) nextState=ch62;
else nextState=ch63;


ch13:if (channel ==6'b001101) nextState=ch13;
else if (channel ==6'b000001) nextState=ch1;
else if (channel ==6'b000010) nextState=ch2;
else if (channel ==6'b000011) nextState=ch3;
else if (channel ==6'b000100) nextState=ch4;
else if (channel ==6'b000101) nextState=ch5;
else if (channel ==6'b000110) nextState=ch6;
else if (channel ==6'b000111) nextState=ch7;
else if (channel ==6'b001000) nextState=ch8;
else if (channel ==6'b001001) nextState=ch9;
else if (channel ==6'b001010) nextState=ch10;
else if (channel ==6'b001011) nextState=ch11;
else if (channel ==6'b001100) nextState=ch12;
else if (channel ==6'b000000) nextState=ch0;
else if (channel ==6'b001110) nextState=ch14;
else if (channel ==6'b001111) nextState=ch15;
else if (channel ==6'b010000) nextState=ch16;
else if (channel ==6'b010001) nextState=ch17;
else if (channel ==6'b010010) nextState=ch18;
else if (channel ==6'b010011) nextState=ch19;
else if (channel ==6'b010100) nextState=ch20;
else if (channel ==6'b010101) nextState=ch21;
else if (channel ==6'b010110) nextState=ch22;
else if (channel ==6'b010111) nextState=ch23;
else if (channel ==6'b011000) nextState=ch24;
else if (channel ==6'b011001) nextState=ch25;
else if (channel ==6'b011010) nextState=ch26;
else if (channel ==6'b011011) nextState=ch27;
else if (channel ==6'b011100) nextState=ch28;
else if (channel ==6'b011101) nextState=ch29;
else if (channel ==6'b011110) nextState=ch30;
else if (channel ==6'b011111) nextState=ch31;
else if (channel ==6'b100000) nextState=ch32;
else if (channel ==6'b100001) nextState=ch33;
else if (channel ==6'b100010) nextState=ch34;
else if (channel ==6'b100011) nextState=ch35;
else if (channel ==6'b100100) nextState=ch36;
else if (channel ==6'b100101) nextState=ch37;
else if (channel ==6'b100110) nextState=ch38;
else if (channel ==6'b100111) nextState=ch39;
else if (channel ==6'b101000) nextState=ch40;
else if (channel ==6'b101001) nextState=ch41;
else if (channel ==6'b101010) nextState=ch42;
else if (channel ==6'b101011) nextState=ch43;
else if (channel ==6'b101100) nextState=ch44;
else if (channel ==6'b101101) nextState=ch45;
else if (channel ==6'b101110) nextState=ch46;
else if (channel ==6'b101111) nextState=ch47;
else if (channel ==6'b110000) nextState=ch48;
else if (channel ==6'b110001) nextState=ch49;
else if (channel ==6'b110010) nextState=ch50;
else if (channel ==6'b110011) nextState=ch51;
else if (channel ==6'b110100) nextState=ch52;
else if (channel ==6'b110101) nextState=ch53;
else if (channel ==6'b110110) nextState=ch54;
else if (channel ==6'b110111) nextState=ch55;
else if (channel ==6'b111000) nextState=ch56;
else if (channel ==6'b111001) nextState=ch57;
else if (channel ==6'b111010) nextState=ch58;
else if (channel ==6'b111011) nextState=ch59;
else if (channel ==6'b111100) nextState=ch60;
else if (channel ==6'b111101) nextState=ch61;
else if (channel ==6'b111110) nextState=ch62;
else nextState=ch63;


ch14:if (channel ==6'b001110) nextState=ch14;
else if (channel ==6'b000001) nextState=ch1;
else if (channel ==6'b000010) nextState=ch2;
else if (channel ==6'b000011) nextState=ch3;
else if (channel ==6'b000100) nextState=ch4;
else if (channel ==6'b000101) nextState=ch5;
else if (channel ==6'b000110) nextState=ch6;
else if (channel ==6'b000111) nextState=ch7;
else if (channel ==6'b001000) nextState=ch8;
else if (channel ==6'b001001) nextState=ch9;
else if (channel ==6'b001010) nextState=ch10;
else if (channel ==6'b001011) nextState=ch11;
else if (channel ==6'b001100) nextState=ch12;
else if (channel ==6'b001101) nextState=ch13;
else if (channel ==6'b000000) nextState=ch0;
else if (channel ==6'b001111) nextState=ch15;
else if (channel ==6'b010000) nextState=ch16;
else if (channel ==6'b010001) nextState=ch17;
else if (channel ==6'b010010) nextState=ch18;
else if (channel ==6'b010011) nextState=ch19;
else if (channel ==6'b010100) nextState=ch20;
else if (channel ==6'b010101) nextState=ch21;
else if (channel ==6'b010110) nextState=ch22;
else if (channel ==6'b010111) nextState=ch23;
else if (channel ==6'b011000) nextState=ch24;
else if (channel ==6'b011001) nextState=ch25;
else if (channel ==6'b011010) nextState=ch26;
else if (channel ==6'b011011) nextState=ch27;
else if (channel ==6'b011100) nextState=ch28;
else if (channel ==6'b011101) nextState=ch29;
else if (channel ==6'b011110) nextState=ch30;
else if (channel ==6'b011111) nextState=ch31;
else if (channel ==6'b100000) nextState=ch32;
else if (channel ==6'b100001) nextState=ch33;
else if (channel ==6'b100010) nextState=ch34;
else if (channel ==6'b100011) nextState=ch35;
else if (channel ==6'b100100) nextState=ch36;
else if (channel ==6'b100101) nextState=ch37;
else if (channel ==6'b100110) nextState=ch38;
else if (channel ==6'b100111) nextState=ch39;
else if (channel ==6'b101000) nextState=ch40;
else if (channel ==6'b101001) nextState=ch41;
else if (channel ==6'b101010) nextState=ch42;
else if (channel ==6'b101011) nextState=ch43;
else if (channel ==6'b101100) nextState=ch44;
else if (channel ==6'b101101) nextState=ch45;
else if (channel ==6'b101110) nextState=ch46;
else if (channel ==6'b101111) nextState=ch47;
else if (channel ==6'b110000) nextState=ch48;
else if (channel ==6'b110001) nextState=ch49;
else if (channel ==6'b110010) nextState=ch50;
else if (channel ==6'b110011) nextState=ch51;
else if (channel ==6'b110100) nextState=ch52;
else if (channel ==6'b110101) nextState=ch53;
else if (channel ==6'b110110) nextState=ch54;
else if (channel ==6'b110111) nextState=ch55;
else if (channel ==6'b111000) nextState=ch56;
else if (channel ==6'b111001) nextState=ch57;
else if (channel ==6'b111010) nextState=ch58;
else if (channel ==6'b111011) nextState=ch59;
else if (channel ==6'b111100) nextState=ch60;
else if (channel ==6'b111101) nextState=ch61;
else if (channel ==6'b111110) nextState=ch62;
else nextState=ch63;


ch15:if (channel==6'b001111) nextState=ch15;
else if (channel ==6'b000001) nextState=ch1;
else if (channel ==6'b000010) nextState=ch2;
else if (channel ==6'b000011) nextState=ch3;
else if (channel ==6'b000100) nextState=ch4;
else if (channel ==6'b000101) nextState=ch5;
else if (channel ==6'b000110) nextState=ch6;
else if (channel ==6'b000111) nextState=ch7;
else if (channel ==6'b001000) nextState=ch8;
else if (channel ==6'b001001) nextState=ch9;
else if (channel ==6'b001010) nextState=ch10;
else if (channel ==6'b001011) nextState=ch11;
else if (channel ==6'b001100) nextState=ch12;
else if (channel ==6'b001101) nextState=ch13;
else if (channel ==6'b001110) nextState=ch14;
else if (channel ==6'b000000) nextState=ch0;
else if (channel ==6'b010000) nextState=ch16;
else if (channel ==6'b010001) nextState=ch17;
else if (channel ==6'b010010) nextState=ch18;
else if (channel ==6'b010011) nextState=ch19;
else if (channel ==6'b010100) nextState=ch20;
else if (channel ==6'b010101) nextState=ch21;
else if (channel ==6'b010110) nextState=ch22;
else if (channel ==6'b010111) nextState=ch23;
else if (channel ==6'b011000) nextState=ch24;
else if (channel ==6'b011001) nextState=ch25;
else if (channel ==6'b011010) nextState=ch26;
else if (channel ==6'b011011) nextState=ch27;
else if (channel ==6'b011100) nextState=ch28;
else if (channel ==6'b011101) nextState=ch29;
else if (channel ==6'b011110) nextState=ch30;
else if (channel ==6'b011111) nextState=ch31;
else if (channel ==6'b100000) nextState=ch32;
else if (channel ==6'b100001) nextState=ch33;
else if (channel ==6'b100010) nextState=ch34;
else if (channel ==6'b100011) nextState=ch35;
else if (channel ==6'b100100) nextState=ch36;
else if (channel ==6'b100101) nextState=ch37;
else if (channel ==6'b100110) nextState=ch38;
else if (channel ==6'b100111) nextState=ch39;
else if (channel ==6'b101000) nextState=ch40;
else if (channel ==6'b101001) nextState=ch41;
else if (channel ==6'b101010) nextState=ch42;
else if (channel ==6'b101011) nextState=ch43;
else if (channel ==6'b101100) nextState=ch44;
else if (channel ==6'b101101) nextState=ch45;
else if (channel ==6'b101110) nextState=ch46;
else if (channel ==6'b101111) nextState=ch47;
else if (channel ==6'b110000) nextState=ch48;
else if (channel ==6'b110001) nextState=ch49;
else if (channel ==6'b110010) nextState=ch50;
else if (channel ==6'b110011) nextState=ch51;
else if (channel ==6'b110100) nextState=ch52;
else if (channel ==6'b110101) nextState=ch53;
else if (channel ==6'b110110) nextState=ch54;
else if (channel ==6'b110111) nextState=ch55;
else if (channel ==6'b111000) nextState=ch56;
else if (channel ==6'b111001) nextState=ch57;
else if (channel ==6'b111010) nextState=ch58;
else if (channel ==6'b111011) nextState=ch59;
else if (channel ==6'b111100) nextState=ch60;
else if (channel ==6'b111101) nextState=ch61;
else if (channel ==6'b111110) nextState=ch62;
else nextState=ch63;


ch16:if (channel ==6'b010000) nextState=ch16;
else if (channel ==6'b000001) nextState=ch1;
else if (channel ==6'b000010) nextState=ch2;
else if (channel ==6'b000011) nextState=ch3;
else if (channel ==6'b000100) nextState=ch4;
else if (channel ==6'b000101) nextState=ch5;
else if (channel ==6'b000110) nextState=ch6;
else if (channel ==6'b000111) nextState=ch7;
else if (channel ==6'b001000) nextState=ch8;
else if (channel ==6'b001001) nextState=ch9;
else if (channel ==6'b001010) nextState=ch10;
else if (channel ==6'b001011) nextState=ch11;
else if (channel ==6'b001100) nextState=ch12;
else if (channel ==6'b001101) nextState=ch13;
else if (channel ==6'b001110) nextState=ch14;
else if (channel ==6'b001111) nextState=ch15;
else if (channel ==6'b000000) nextState=ch0;
else if (channel ==6'b010001) nextState=ch17;
else if (channel ==6'b010010) nextState=ch18;
else if (channel ==6'b010011) nextState=ch19;
else if (channel ==6'b010100) nextState=ch20;
else if (channel ==6'b010101) nextState=ch21;
else if (channel ==6'b010110) nextState=ch22;
else if (channel ==6'b010111) nextState=ch23;
else if (channel ==6'b011000) nextState=ch24;
else if (channel ==6'b011001) nextState=ch25;
else if (channel ==6'b011010) nextState=ch26;
else if (channel ==6'b011011) nextState=ch27;
else if (channel ==6'b011100) nextState=ch28;
else if (channel ==6'b011101) nextState=ch29;
else if (channel ==6'b011110) nextState=ch30;
else if (channel ==6'b011111) nextState=ch31;
else if (channel ==6'b100000) nextState=ch32;
else if (channel ==6'b100001) nextState=ch33;
else if (channel ==6'b100010) nextState=ch34;
else if (channel ==6'b100011) nextState=ch35;
else if (channel ==6'b100100) nextState=ch36;
else if (channel ==6'b100101) nextState=ch37;
else if (channel ==6'b100110) nextState=ch38;
else if (channel ==6'b100111) nextState=ch39;
else if (channel ==6'b101000) nextState=ch40;
else if (channel ==6'b101001) nextState=ch41;
else if (channel ==6'b101010) nextState=ch42;
else if (channel ==6'b101011) nextState=ch43;
else if (channel ==6'b101100) nextState=ch44;
else if (channel ==6'b101101) nextState=ch45;
else if (channel ==6'b101110) nextState=ch46;
else if (channel ==6'b101111) nextState=ch47;
else if (channel ==6'b110000) nextState=ch48;
else if (channel ==6'b110001) nextState=ch49;
else if (channel ==6'b110010) nextState=ch50;
else if (channel ==6'b110011) nextState=ch51;
else if (channel ==6'b110100) nextState=ch52;
else if (channel ==6'b110101) nextState=ch53;
else if (channel ==6'b110110) nextState=ch54;
else if (channel ==6'b110111) nextState=ch55;
else if (channel ==6'b111000) nextState=ch56;
else if (channel ==6'b111001) nextState=ch57;
else if (channel ==6'b111010) nextState=ch58;
else if (channel ==6'b111011) nextState=ch59;
else if (channel ==6'b111100) nextState=ch60;
else if (channel ==6'b111101) nextState=ch61;
else if (channel ==6'b111110) nextState=ch62;
else nextState=ch63;


ch17:if (channel ==6'b010001) nextState=ch17;
else if (channel ==6'b000001) nextState=ch1;
else if (channel ==6'b000010) nextState=ch2;
else if (channel ==6'b000011) nextState=ch3;
else if (channel ==6'b000100) nextState=ch4;
else if (channel ==6'b000101) nextState=ch5;
else if (channel ==6'b000110) nextState=ch6;
else if (channel ==6'b000111) nextState=ch7;
else if (channel ==6'b001000) nextState=ch8;
else if (channel ==6'b001001) nextState=ch9;
else if (channel ==6'b001010) nextState=ch10;
else if (channel ==6'b001011) nextState=ch11;
else if (channel ==6'b001100) nextState=ch12;
else if (channel ==6'b001101) nextState=ch13;
else if (channel ==6'b001110) nextState=ch14;
else if (channel ==6'b001111) nextState=ch15;
else if (channel ==6'b010000) nextState=ch16;
else if (channel ==6'b000000) nextState=ch0;
else if (channel ==6'b010010) nextState=ch18;
else if (channel ==6'b010011) nextState=ch19;
else if (channel ==6'b010100) nextState=ch20;
else if (channel ==6'b010101) nextState=ch21;
else if (channel ==6'b010110) nextState=ch22;
else if (channel ==6'b010111) nextState=ch23;
else if (channel ==6'b011000) nextState=ch24;
else if (channel ==6'b011001) nextState=ch25;
else if (channel ==6'b011010) nextState=ch26;
else if (channel ==6'b011011) nextState=ch27;
else if (channel ==6'b011100) nextState=ch28;
else if (channel ==6'b011101) nextState=ch29;
else if (channel ==6'b011110) nextState=ch30;
else if (channel ==6'b011111) nextState=ch31;
else if (channel ==6'b100000) nextState=ch32;
else if (channel ==6'b100001) nextState=ch33;
else if (channel ==6'b100010) nextState=ch34;
else if (channel ==6'b100011) nextState=ch35;
else if (channel ==6'b100100) nextState=ch36;
else if (channel ==6'b100101) nextState=ch37;
else if (channel ==6'b100110) nextState=ch38;
else if (channel ==6'b100111) nextState=ch39;
else if (channel ==6'b101000) nextState=ch40;
else if (channel ==6'b101001) nextState=ch41;
else if (channel ==6'b101010) nextState=ch42;
else if (channel ==6'b101011) nextState=ch43;
else if (channel ==6'b101100) nextState=ch44;
else if (channel ==6'b101101) nextState=ch45;
else if (channel ==6'b101110) nextState=ch46;
else if (channel ==6'b101111) nextState=ch47;
else if (channel ==6'b110000) nextState=ch48;
else if (channel ==6'b110001) nextState=ch49;
else if (channel ==6'b110010) nextState=ch50;
else if (channel ==6'b110011) nextState=ch51;
else if (channel ==6'b110100) nextState=ch52;
else if (channel ==6'b110101) nextState=ch53;
else if (channel ==6'b110110) nextState=ch54;
else if (channel ==6'b110111) nextState=ch55;
else if (channel ==6'b111000) nextState=ch56;
else if (channel ==6'b111001) nextState=ch57;
else if (channel ==6'b111010) nextState=ch58;
else if (channel ==6'b111011) nextState=ch59;
else if (channel ==6'b111100) nextState=ch60;
else if (channel ==6'b111101) nextState=ch61;
else if (channel ==6'b111110) nextState=ch62;
else nextState=ch63;


ch18:if (channel ==6'b010010) nextState=ch18;
else if (channel ==6'b000001) nextState=ch1;
else if (channel ==6'b000010) nextState=ch2;
else if (channel ==6'b000011) nextState=ch3;
else if (channel ==6'b000100) nextState=ch4;
else if (channel ==6'b000101) nextState=ch5;
else if (channel ==6'b000110) nextState=ch6;
else if (channel ==6'b000111) nextState=ch7;
else if (channel ==6'b001000) nextState=ch8;
else if (channel ==6'b001001) nextState=ch9;
else if (channel ==6'b001010) nextState=ch10;
else if (channel ==6'b001011) nextState=ch11;
else if (channel ==6'b001100) nextState=ch12;
else if (channel ==6'b001101) nextState=ch13;
else if (channel ==6'b001110) nextState=ch14;
else if (channel ==6'b001111) nextState=ch15;
else if (channel ==6'b010000) nextState=ch16;
else if (channel ==6'b010001) nextState=ch17;
else if (channel ==6'b000000) nextState=ch0;
else if (channel ==6'b010011) nextState=ch19;
else if (channel ==6'b010100) nextState=ch20;
else if (channel ==6'b010101) nextState=ch21;
else if (channel ==6'b010110) nextState=ch22;
else if (channel ==6'b010111) nextState=ch23;
else if (channel ==6'b011000) nextState=ch24;
else if (channel ==6'b011001) nextState=ch25;
else if (channel ==6'b011010) nextState=ch26;
else if (channel ==6'b011011) nextState=ch27;
else if (channel ==6'b011100) nextState=ch28;
else if (channel ==6'b011101) nextState=ch29;
else if (channel ==6'b011110) nextState=ch30;
else if (channel ==6'b011111) nextState=ch31;
else if (channel ==6'b100000) nextState=ch32;
else if (channel ==6'b100001) nextState=ch33;
else if (channel ==6'b100010) nextState=ch34;
else if (channel ==6'b100011) nextState=ch35;
else if (channel ==6'b100100) nextState=ch36;
else if (channel ==6'b100101) nextState=ch37;
else if (channel ==6'b100110) nextState=ch38;
else if (channel ==6'b100111) nextState=ch39;
else if (channel ==6'b101000) nextState=ch40;
else if (channel ==6'b101001) nextState=ch41;
else if (channel ==6'b101010) nextState=ch42;
else if (channel ==6'b101011) nextState=ch43;
else if (channel ==6'b101100) nextState=ch44;
else if (channel ==6'b101101) nextState=ch45;
else if (channel ==6'b101110) nextState=ch46;
else if (channel ==6'b101111) nextState=ch47;
else if (channel ==6'b110000) nextState=ch48;
else if (channel ==6'b110001) nextState=ch49;
else if (channel ==6'b110010) nextState=ch50;
else if (channel ==6'b110011) nextState=ch51;
else if (channel ==6'b110100) nextState=ch52;
else if (channel ==6'b110101) nextState=ch53;
else if (channel ==6'b110110) nextState=ch54;
else if (channel ==6'b110111) nextState=ch55;
else if (channel ==6'b111000) nextState=ch56;
else if (channel ==6'b111001) nextState=ch57;
else if (channel ==6'b111010) nextState=ch58;
else if (channel ==6'b111011) nextState=ch59;
else if (channel ==6'b111100) nextState=ch60;
else if (channel ==6'b111101) nextState=ch61;
else if (channel ==6'b111110) nextState=ch62;
else nextState=ch63;


ch19:if (channel ==6'b010011) nextState=ch19;
else if (channel ==6'b000001) nextState=ch1;
else if (channel ==6'b000010) nextState=ch2;
else if (channel ==6'b000011) nextState=ch3;
else if (channel ==6'b000100) nextState=ch4;
else if (channel ==6'b000101) nextState=ch5;
else if (channel ==6'b000110) nextState=ch6;
else if (channel ==6'b000111) nextState=ch7;
else if (channel ==6'b001000) nextState=ch8;
else if (channel ==6'b001001) nextState=ch9;
else if (channel ==6'b001010) nextState=ch10;
else if (channel ==6'b001011) nextState=ch11;
else if (channel ==6'b001100) nextState=ch12;
else if (channel ==6'b001101) nextState=ch13;
else if (channel ==6'b001110) nextState=ch14;
else if (channel ==6'b001111) nextState=ch15;
else if (channel ==6'b010000) nextState=ch16;
else if (channel ==6'b010001) nextState=ch17;
else if (channel ==6'b010010) nextState=ch18;
else if (channel ==6'b000000) nextState=ch0;
else if (channel ==6'b010100) nextState=ch20;
else if (channel ==6'b010101) nextState=ch21;
else if (channel ==6'b010110) nextState=ch22;
else if (channel ==6'b010111) nextState=ch23;
else if (channel ==6'b011000) nextState=ch24;
else if (channel ==6'b011001) nextState=ch25;
else if (channel ==6'b011010) nextState=ch26;
else if (channel ==6'b011011) nextState=ch27;
else if (channel ==6'b011100) nextState=ch28;
else if (channel ==6'b011101) nextState=ch29;
else if (channel ==6'b011110) nextState=ch30;
else if (channel ==6'b011111) nextState=ch31;
else if (channel ==6'b100000) nextState=ch32;
else if (channel ==6'b100001) nextState=ch33;
else if (channel ==6'b100010) nextState=ch34;
else if (channel ==6'b100011) nextState=ch35;
else if (channel ==6'b100100) nextState=ch36;
else if (channel ==6'b100101) nextState=ch37;
else if (channel ==6'b100110) nextState=ch38;
else if (channel ==6'b100111) nextState=ch39;
else if (channel ==6'b101000) nextState=ch40;
else if (channel ==6'b101001) nextState=ch41;
else if (channel ==6'b101010) nextState=ch42;
else if (channel ==6'b101011) nextState=ch43;
else if (channel ==6'b101100) nextState=ch44;
else if (channel ==6'b101101) nextState=ch45;
else if (channel ==6'b101110) nextState=ch46;
else if (channel ==6'b101111) nextState=ch47;
else if (channel ==6'b110000) nextState=ch48;
else if (channel ==6'b110001) nextState=ch49;
else if (channel ==6'b110010) nextState=ch50;
else if (channel ==6'b110011) nextState=ch51;
else if (channel ==6'b110100) nextState=ch52;
else if (channel ==6'b110101) nextState=ch53;
else if (channel ==6'b110110) nextState=ch54;
else if (channel ==6'b110111) nextState=ch55;
else if (channel ==6'b111000) nextState=ch56;
else if (channel ==6'b111001) nextState=ch57;
else if (channel ==6'b111010) nextState=ch58;
else if (channel ==6'b111011) nextState=ch59;
else if (channel ==6'b111100) nextState=ch60;
else if (channel ==6'b111101) nextState=ch61;
else if (channel ==6'b111110) nextState=ch62;
else nextState=ch63;


ch20:if (channel ==6'b010100) nextState=ch20;
else if (channel ==6'b000001) nextState=ch1;
else if (channel ==6'b000010) nextState=ch2;
else if (channel ==6'b000011) nextState=ch3;
else if (channel ==6'b000100) nextState=ch4;
else if (channel ==6'b000101) nextState=ch5;
else if (channel ==6'b000110) nextState=ch6;
else if (channel ==6'b000111) nextState=ch7;
else if (channel ==6'b001000) nextState=ch8;
else if (channel ==6'b001001) nextState=ch9;
else if (channel ==6'b001010) nextState=ch10;
else if (channel ==6'b001011) nextState=ch11;
else if (channel ==6'b001100) nextState=ch12;
else if (channel ==6'b001101) nextState=ch13;
else if (channel ==6'b001110) nextState=ch14;
else if (channel ==6'b001111) nextState=ch15;
else if (channel ==6'b010000) nextState=ch16;
else if (channel ==6'b010001) nextState=ch17;
else if (channel ==6'b010010) nextState=ch18;
else if (channel ==6'b010011) nextState=ch19;
else if (channel ==6'b000000) nextState=ch0;
else if (channel ==6'b010101) nextState=ch21;
else if (channel ==6'b010110) nextState=ch22;
else if (channel ==6'b010111) nextState=ch23;
else if (channel ==6'b011000) nextState=ch24;
else if (channel ==6'b011001) nextState=ch25;
else if (channel ==6'b011010) nextState=ch26;
else if (channel ==6'b011011) nextState=ch27;
else if (channel ==6'b011100) nextState=ch28;
else if (channel ==6'b011101) nextState=ch29;
else if (channel ==6'b011110) nextState=ch30;
else if (channel ==6'b011111) nextState=ch31;
else if (channel ==6'b100000) nextState=ch32;
else if (channel ==6'b100001) nextState=ch33;
else if (channel ==6'b100010) nextState=ch34;
else if (channel ==6'b100011) nextState=ch35;
else if (channel ==6'b100100) nextState=ch36;
else if (channel ==6'b100101) nextState=ch37;
else if (channel ==6'b100110) nextState=ch38;
else if (channel ==6'b100111) nextState=ch39;
else if (channel ==6'b101000) nextState=ch40;
else if (channel ==6'b101001) nextState=ch41;
else if (channel ==6'b101010) nextState=ch42;
else if (channel ==6'b101011) nextState=ch43;
else if (channel ==6'b101100) nextState=ch44;
else if (channel ==6'b101101) nextState=ch45;
else if (channel ==6'b101110) nextState=ch46;
else if (channel ==6'b101111) nextState=ch47;
else if (channel ==6'b110000) nextState=ch48;
else if (channel ==6'b110001) nextState=ch49;
else if (channel ==6'b110010) nextState=ch50;
else if (channel ==6'b110011) nextState=ch51;
else if (channel ==6'b110100) nextState=ch52;
else if (channel ==6'b110101) nextState=ch53;
else if (channel ==6'b110110) nextState=ch54;
else if (channel ==6'b110111) nextState=ch55;
else if (channel ==6'b111000) nextState=ch56;
else if (channel ==6'b111001) nextState=ch57;
else if (channel ==6'b111010) nextState=ch58;
else if (channel ==6'b111011) nextState=ch59;
else if (channel ==6'b111100) nextState=ch60;
else if (channel ==6'b111101) nextState=ch61;
else if (channel ==6'b111110) nextState=ch62;
else nextState=ch63;


ch21:if (channel ==6'b010101) nextState=ch21;
else if (channel ==6'b000001) nextState=ch1;
else if (channel ==6'b000010) nextState=ch2;
else if (channel ==6'b000011) nextState=ch3;
else if (channel ==6'b000100) nextState=ch4;
else if (channel ==6'b000101) nextState=ch5;
else if (channel ==6'b000110) nextState=ch6;
else if (channel ==6'b000111) nextState=ch7;
else if (channel ==6'b001000) nextState=ch8;
else if (channel ==6'b001001) nextState=ch9;
else if (channel ==6'b001010) nextState=ch10;
else if (channel ==6'b001011) nextState=ch11;
else if (channel ==6'b001100) nextState=ch12;
else if (channel ==6'b001101) nextState=ch13;
else if (channel ==6'b001110) nextState=ch14;
else if (channel ==6'b001111) nextState=ch15;
else if (channel ==6'b010000) nextState=ch16;
else if (channel ==6'b010001) nextState=ch17;
else if (channel ==6'b010010) nextState=ch18;
else if (channel ==6'b010011) nextState=ch19;
else if (channel ==6'b010100) nextState=ch20;
else if (channel ==6'b000000) nextState=ch0;
else if (channel ==6'b010110) nextState=ch22;
else if (channel ==6'b010111) nextState=ch23;
else if (channel ==6'b011000) nextState=ch24;
else if (channel ==6'b011001) nextState=ch25;
else if (channel ==6'b011010) nextState=ch26;
else if (channel ==6'b011011) nextState=ch27;
else if (channel ==6'b011100) nextState=ch28;
else if (channel ==6'b011101) nextState=ch29;
else if (channel ==6'b011110) nextState=ch30;
else if (channel ==6'b011111) nextState=ch31;
else if (channel ==6'b100000) nextState=ch32;
else if (channel ==6'b100001) nextState=ch33;
else if (channel ==6'b100010) nextState=ch34;
else if (channel ==6'b100011) nextState=ch35;
else if (channel ==6'b100100) nextState=ch36;
else if (channel ==6'b100101) nextState=ch37;
else if (channel ==6'b100110) nextState=ch38;
else if (channel ==6'b100111) nextState=ch39;
else if (channel ==6'b101000) nextState=ch40;
else if (channel ==6'b101001) nextState=ch41;
else if (channel ==6'b101010) nextState=ch42;
else if (channel ==6'b101011) nextState=ch43;
else if (channel ==6'b101100) nextState=ch44;
else if (channel ==6'b101101) nextState=ch45;
else if (channel ==6'b101110) nextState=ch46;
else if (channel ==6'b101111) nextState=ch47;
else if (channel ==6'b110000) nextState=ch48;
else if (channel ==6'b110001) nextState=ch49;
else if (channel ==6'b110010) nextState=ch50;
else if (channel ==6'b110011) nextState=ch51;
else if (channel ==6'b110100) nextState=ch52;
else if (channel ==6'b110101) nextState=ch53;
else if (channel ==6'b110110) nextState=ch54;
else if (channel ==6'b110111) nextState=ch55;
else if (channel ==6'b111000) nextState=ch56;
else if (channel ==6'b111001) nextState=ch57;
else if (channel ==6'b111010) nextState=ch58;
else if (channel ==6'b111011) nextState=ch59;
else if (channel ==6'b111100) nextState=ch60;
else if (channel ==6'b111101) nextState=ch61;
else if (channel ==6'b111110) nextState=ch62;
else nextState=ch63;


ch22:if (channel ==6'b010110) nextState=ch22;
else if (channel ==6'b000001) nextState=ch1;
else if (channel ==6'b000010) nextState=ch2;
else if (channel ==6'b000011) nextState=ch3;
else if (channel ==6'b000100) nextState=ch4;
else if (channel ==6'b000101) nextState=ch5;
else if (channel ==6'b000110) nextState=ch6;
else if (channel ==6'b000111) nextState=ch7;
else if (channel ==6'b001000) nextState=ch8;
else if (channel ==6'b001001) nextState=ch9;
else if (channel ==6'b001010) nextState=ch10;
else if (channel ==6'b001011) nextState=ch11;
else if (channel ==6'b001100) nextState=ch12;
else if (channel ==6'b001101) nextState=ch13;
else if (channel ==6'b001110) nextState=ch14;
else if (channel ==6'b001111) nextState=ch15;
else if (channel ==6'b010000) nextState=ch16;
else if (channel ==6'b010001) nextState=ch17;
else if (channel ==6'b010010) nextState=ch18;
else if (channel ==6'b010011) nextState=ch19;
else if (channel ==6'b010100) nextState=ch20;
else if (channel ==6'b010101) nextState=ch21;
else if (channel ==6'b000000) nextState=ch0;
else if (channel ==6'b010111) nextState=ch23;
else if (channel ==6'b011000) nextState=ch24;
else if (channel ==6'b011001) nextState=ch25;
else if (channel ==6'b011010) nextState=ch26;
else if (channel ==6'b011011) nextState=ch27;
else if (channel ==6'b011100) nextState=ch28;
else if (channel ==6'b011101) nextState=ch29;
else if (channel ==6'b011110) nextState=ch30;
else if (channel ==6'b011111) nextState=ch31;
else if (channel ==6'b100000) nextState=ch32;
else if (channel ==6'b100001) nextState=ch33;
else if (channel ==6'b100010) nextState=ch34;
else if (channel ==6'b100011) nextState=ch35;
else if (channel ==6'b100100) nextState=ch36;
else if (channel ==6'b100101) nextState=ch37;
else if (channel ==6'b100110) nextState=ch38;
else if (channel ==6'b100111) nextState=ch39;
else if (channel ==6'b101000) nextState=ch40;
else if (channel ==6'b101001) nextState=ch41;
else if (channel ==6'b101010) nextState=ch42;
else if (channel ==6'b101011) nextState=ch43;
else if (channel ==6'b101100) nextState=ch44;
else if (channel ==6'b101101) nextState=ch45;
else if (channel ==6'b101110) nextState=ch46;
else if (channel ==6'b101111) nextState=ch47;
else if (channel ==6'b110000) nextState=ch48;
else if (channel ==6'b110001) nextState=ch49;
else if (channel ==6'b110010) nextState=ch50;
else if (channel ==6'b110011) nextState=ch51;
else if (channel ==6'b110100) nextState=ch52;
else if (channel ==6'b110101) nextState=ch53;
else if (channel ==6'b110110) nextState=ch54;
else if (channel ==6'b110111) nextState=ch55;
else if (channel ==6'b111000) nextState=ch56;
else if (channel ==6'b111001) nextState=ch57;
else if (channel ==6'b111010) nextState=ch58;
else if (channel ==6'b111011) nextState=ch59;
else if (channel ==6'b111100) nextState=ch60;
else if (channel ==6'b111101) nextState=ch61;
else if (channel ==6'b111110) nextState=ch62;
else nextState=ch63;


ch23:if (channel ==6'b010111) nextState=ch23;
else if (channel ==6'b000001) nextState=ch1;
else if (channel ==6'b000010) nextState=ch2;
else if (channel ==6'b000011) nextState=ch3;
else if (channel ==6'b000100) nextState=ch4;
else if (channel ==6'b000101) nextState=ch5;
else if (channel ==6'b000110) nextState=ch6;
else if (channel ==6'b000111) nextState=ch7;
else if (channel ==6'b001000) nextState=ch8;
else if (channel ==6'b001001) nextState=ch9;
else if (channel ==6'b001010) nextState=ch10;
else if (channel ==6'b001011) nextState=ch11;
else if (channel ==6'b001100) nextState=ch12;
else if (channel ==6'b001101) nextState=ch13;
else if (channel ==6'b001110) nextState=ch14;
else if (channel ==6'b001111) nextState=ch15;
else if (channel ==6'b010000) nextState=ch16;
else if (channel ==6'b010001) nextState=ch17;
else if (channel ==6'b010010) nextState=ch18;
else if (channel ==6'b010011) nextState=ch19;
else if (channel ==6'b010100) nextState=ch20;
else if (channel ==6'b010101) nextState=ch21;
else if (channel ==6'b010110) nextState=ch22;
else if (channel ==6'b000000) nextState=ch0;
else if (channel ==6'b011000) nextState=ch24;
else if (channel ==6'b011001) nextState=ch25;
else if (channel ==6'b011010) nextState=ch26;
else if (channel ==6'b011011) nextState=ch27;
else if (channel ==6'b011100) nextState=ch28;
else if (channel ==6'b011101) nextState=ch29;
else if (channel ==6'b011110) nextState=ch30;
else if (channel ==6'b011111) nextState=ch31;
else if (channel ==6'b100000) nextState=ch32;
else if (channel ==6'b100001) nextState=ch33;
else if (channel ==6'b100010) nextState=ch34;
else if (channel ==6'b100011) nextState=ch35;
else if (channel ==6'b100100) nextState=ch36;
else if (channel ==6'b100101) nextState=ch37;
else if (channel ==6'b100110) nextState=ch38;
else if (channel ==6'b100111) nextState=ch39;
else if (channel ==6'b101000) nextState=ch40;
else if (channel ==6'b101001) nextState=ch41;
else if (channel ==6'b101010) nextState=ch42;
else if (channel ==6'b101011) nextState=ch43;
else if (channel ==6'b101100) nextState=ch44;
else if (channel ==6'b101101) nextState=ch45;
else if (channel ==6'b101110) nextState=ch46;
else if (channel ==6'b101111) nextState=ch47;
else if (channel ==6'b110000) nextState=ch48;
else if (channel ==6'b110001) nextState=ch49;
else if (channel ==6'b110010) nextState=ch50;
else if (channel ==6'b110011) nextState=ch51;
else if (channel ==6'b110100) nextState=ch52;
else if (channel ==6'b110101) nextState=ch53;
else if (channel ==6'b110110) nextState=ch54;
else if (channel ==6'b110111) nextState=ch55;
else if (channel ==6'b111000) nextState=ch56;
else if (channel ==6'b111001) nextState=ch57;
else if (channel ==6'b111010) nextState=ch58;
else if (channel ==6'b111011) nextState=ch59;
else if (channel ==6'b111100) nextState=ch60;
else if (channel ==6'b111101) nextState=ch61;
else if (channel ==6'b111110) nextState=ch62;
else nextState=ch63;


ch24:if (channel ==6'b011000) nextState=ch24;
else if (channel ==6'b000001) nextState=ch1;
else if (channel ==6'b000010) nextState=ch2;
else if (channel ==6'b000011) nextState=ch3;
else if (channel ==6'b000100) nextState=ch4;
else if (channel ==6'b000101) nextState=ch5;
else if (channel ==6'b000110) nextState=ch6;
else if (channel ==6'b000111) nextState=ch7;
else if (channel ==6'b001000) nextState=ch8;
else if (channel ==6'b001001) nextState=ch9;
else if (channel ==6'b001010) nextState=ch10;
else if (channel ==6'b001011) nextState=ch11;
else if (channel ==6'b001100) nextState=ch12;
else if (channel ==6'b001101) nextState=ch13;
else if (channel ==6'b001110) nextState=ch14;
else if (channel ==6'b001111) nextState=ch15;
else if (channel ==6'b010000) nextState=ch16;
else if (channel ==6'b010001) nextState=ch17;
else if (channel ==6'b010010) nextState=ch18;
else if (channel ==6'b010011) nextState=ch19;
else if (channel ==6'b010100) nextState=ch20;
else if (channel ==6'b010101) nextState=ch21;
else if (channel ==6'b010110) nextState=ch22;
else if (channel ==6'b010111) nextState=ch23;
else if (channel ==6'b000000) nextState=ch0;
else if (channel ==6'b011001) nextState=ch25;
else if (channel ==6'b011010) nextState=ch26;
else if (channel ==6'b011011) nextState=ch27;
else if (channel ==6'b011100) nextState=ch28;
else if (channel ==6'b011101) nextState=ch29;
else if (channel ==6'b011110) nextState=ch30;
else if (channel ==6'b011111) nextState=ch31;
else if (channel ==6'b100000) nextState=ch32;
else if (channel ==6'b100001) nextState=ch33;
else if (channel ==6'b100010) nextState=ch34;
else if (channel ==6'b100011) nextState=ch35;
else if (channel ==6'b100100) nextState=ch36;
else if (channel ==6'b100101) nextState=ch37;
else if (channel ==6'b100110) nextState=ch38;
else if (channel ==6'b100111) nextState=ch39;
else if (channel ==6'b101000) nextState=ch40;
else if (channel ==6'b101001) nextState=ch41;
else if (channel ==6'b101010) nextState=ch42;
else if (channel ==6'b101011) nextState=ch43;
else if (channel ==6'b101100) nextState=ch44;
else if (channel ==6'b101101) nextState=ch45;
else if (channel ==6'b101110) nextState=ch46;
else if (channel ==6'b101111) nextState=ch47;
else if (channel ==6'b110000) nextState=ch48;
else if (channel ==6'b110001) nextState=ch49;
else if (channel ==6'b110010) nextState=ch50;
else if (channel ==6'b110011) nextState=ch51;
else if (channel ==6'b110100) nextState=ch52;
else if (channel ==6'b110101) nextState=ch53;
else if (channel ==6'b110110) nextState=ch54;
else if (channel ==6'b110111) nextState=ch55;
else if (channel ==6'b111000) nextState=ch56;
else if (channel ==6'b111001) nextState=ch57;
else if (channel ==6'b111010) nextState=ch58;
else if (channel ==6'b111011) nextState=ch59;
else if (channel ==6'b111100) nextState=ch60;
else if (channel ==6'b111101) nextState=ch61;
else if (channel ==6'b111110) nextState=ch62;
else nextState=ch63;


ch25:if (channel ==6'b011001) nextState=ch25;
else if (channel ==6'b000001) nextState=ch1;
else if (channel ==6'b000010) nextState=ch2;
else if (channel ==6'b000011) nextState=ch3;
else if (channel ==6'b000100) nextState=ch4;
else if (channel ==6'b000101) nextState=ch5;
else if (channel ==6'b000110) nextState=ch6;
else if (channel ==6'b000111) nextState=ch7;
else if (channel ==6'b001000) nextState=ch8;
else if (channel ==6'b001001) nextState=ch9;
else if (channel ==6'b001010) nextState=ch10;
else if (channel ==6'b001011) nextState=ch11;
else if (channel ==6'b001100) nextState=ch12;
else if (channel ==6'b001101) nextState=ch13;
else if (channel ==6'b001110) nextState=ch14;
else if (channel ==6'b001111) nextState=ch15;
else if (channel ==6'b010000) nextState=ch16;
else if (channel ==6'b010001) nextState=ch17;
else if (channel ==6'b010010) nextState=ch18;
else if (channel ==6'b010011) nextState=ch19;
else if (channel ==6'b010100) nextState=ch20;
else if (channel ==6'b010101) nextState=ch21;
else if (channel ==6'b010110) nextState=ch22;
else if (channel ==6'b010111) nextState=ch23;
else if (channel ==6'b011000) nextState=ch24;
else if (channel ==6'b000000) nextState=ch0;
else if (channel ==6'b011010) nextState=ch26;
else if (channel ==6'b011011) nextState=ch27;
else if (channel ==6'b011100) nextState=ch28;
else if (channel ==6'b011101) nextState=ch29;
else if (channel ==6'b011110) nextState=ch30;
else if (channel ==6'b011111) nextState=ch31;
else if (channel ==6'b100000) nextState=ch32;
else if (channel ==6'b100001) nextState=ch33;
else if (channel ==6'b100010) nextState=ch34;
else if (channel ==6'b100011) nextState=ch35;
else if (channel ==6'b100100) nextState=ch36;
else if (channel ==6'b100101) nextState=ch37;
else if (channel ==6'b100110) nextState=ch38;
else if (channel ==6'b100111) nextState=ch39;
else if (channel ==6'b101000) nextState=ch40;
else if (channel ==6'b101001) nextState=ch41;
else if (channel ==6'b101010) nextState=ch42;
else if (channel ==6'b101011) nextState=ch43;
else if (channel ==6'b101100) nextState=ch44;
else if (channel ==6'b101101) nextState=ch45;
else if (channel ==6'b101110) nextState=ch46;
else if (channel ==6'b101111) nextState=ch47;
else if (channel ==6'b110000) nextState=ch48;
else if (channel ==6'b110001) nextState=ch49;
else if (channel ==6'b110010) nextState=ch50;
else if (channel ==6'b110011) nextState=ch51;
else if (channel ==6'b110100) nextState=ch52;
else if (channel ==6'b110101) nextState=ch53;
else if (channel ==6'b110110) nextState=ch54;
else if (channel ==6'b110111) nextState=ch55;
else if (channel ==6'b111000) nextState=ch56;
else if (channel ==6'b111001) nextState=ch57;
else if (channel ==6'b111010) nextState=ch58;
else if (channel ==6'b111011) nextState=ch59;
else if (channel ==6'b111100) nextState=ch60;
else if (channel ==6'b111101) nextState=ch61;
else if (channel ==6'b111110) nextState=ch62;
else nextState=ch63;


ch26:if (channel ==6'b011010) nextState=ch26;
else if (channel ==6'b000001) nextState=ch1;
else if (channel ==6'b000010) nextState=ch2;
else if (channel ==6'b000011) nextState=ch3;
else if (channel ==6'b000100) nextState=ch4;
else if (channel ==6'b000101) nextState=ch5;
else if (channel ==6'b000110) nextState=ch6;
else if (channel ==6'b000111) nextState=ch7;
else if (channel ==6'b001000) nextState=ch8;
else if (channel ==6'b001001) nextState=ch9;
else if (channel ==6'b001010) nextState=ch10;
else if (channel ==6'b001011) nextState=ch11;
else if (channel ==6'b001100) nextState=ch12;
else if (channel ==6'b001101) nextState=ch13;
else if (channel ==6'b001110) nextState=ch14;
else if (channel ==6'b001111) nextState=ch15;
else if (channel ==6'b010000) nextState=ch16;
else if (channel ==6'b010001) nextState=ch17;
else if (channel ==6'b010010) nextState=ch18;
else if (channel ==6'b010011) nextState=ch19;
else if (channel ==6'b010100) nextState=ch20;
else if (channel ==6'b010101) nextState=ch21;
else if (channel ==6'b010110) nextState=ch22;
else if (channel ==6'b010111) nextState=ch23;
else if (channel ==6'b011000) nextState=ch24;
else if (channel ==6'b011001) nextState=ch25;
else if (channel ==6'b000000) nextState=ch0;
else if (channel ==6'b011011) nextState=ch27;
else if (channel ==6'b011100) nextState=ch28;
else if (channel ==6'b011101) nextState=ch29;
else if (channel ==6'b011110) nextState=ch30;
else if (channel ==6'b011111) nextState=ch31;
else if (channel ==6'b100000) nextState=ch32;
else if (channel ==6'b100001) nextState=ch33;
else if (channel ==6'b100010) nextState=ch34;
else if (channel ==6'b100011) nextState=ch35;
else if (channel ==6'b100100) nextState=ch36;
else if (channel ==6'b100101) nextState=ch37;
else if (channel ==6'b100110) nextState=ch38;
else if (channel ==6'b100111) nextState=ch39;
else if (channel ==6'b101000) nextState=ch40;
else if (channel ==6'b101001) nextState=ch41;
else if (channel ==6'b101010) nextState=ch42;
else if (channel ==6'b101011) nextState=ch43;
else if (channel ==6'b101100) nextState=ch44;
else if (channel ==6'b101101) nextState=ch45;
else if (channel ==6'b101110) nextState=ch46;
else if (channel ==6'b101111) nextState=ch47;
else if (channel ==6'b110000) nextState=ch48;
else if (channel ==6'b110001) nextState=ch49;
else if (channel ==6'b110010) nextState=ch50;
else if (channel ==6'b110011) nextState=ch51;
else if (channel ==6'b110100) nextState=ch52;
else if (channel ==6'b110101) nextState=ch53;
else if (channel ==6'b110110) nextState=ch54;
else if (channel ==6'b110111) nextState=ch55;
else if (channel ==6'b111000) nextState=ch56;
else if (channel ==6'b111001) nextState=ch57;
else if (channel ==6'b111010) nextState=ch58;
else if (channel ==6'b111011) nextState=ch59;
else if (channel ==6'b111100) nextState=ch60;
else if (channel ==6'b111101) nextState=ch61;
else if (channel ==6'b111110) nextState=ch62;
else nextState=ch63;


ch27:if (channel ==6'b011011) nextState=ch27;
else if (channel ==6'b000001) nextState=ch1;
else if (channel ==6'b000010) nextState=ch2;
else if (channel ==6'b000011) nextState=ch3;
else if (channel ==6'b000100) nextState=ch4;
else if (channel ==6'b000101) nextState=ch5;
else if (channel ==6'b000110) nextState=ch6;
else if (channel ==6'b000111) nextState=ch7;
else if (channel ==6'b001000) nextState=ch8;
else if (channel ==6'b001001) nextState=ch9;
else if (channel ==6'b001010) nextState=ch10;
else if (channel ==6'b001011) nextState=ch11;
else if (channel ==6'b001100) nextState=ch12;
else if (channel ==6'b001101) nextState=ch13;
else if (channel ==6'b001110) nextState=ch14;
else if (channel ==6'b001111) nextState=ch15;
else if (channel ==6'b010000) nextState=ch16;
else if (channel ==6'b010001) nextState=ch17;
else if (channel ==6'b010010) nextState=ch18;
else if (channel ==6'b010011) nextState=ch19;
else if (channel ==6'b010100) nextState=ch20;
else if (channel ==6'b010101) nextState=ch21;
else if (channel ==6'b010110) nextState=ch22;
else if (channel ==6'b010111) nextState=ch23;
else if (channel ==6'b011000) nextState=ch24;
else if (channel ==6'b011001) nextState=ch25;
else if (channel ==6'b011010) nextState=ch26;
else if (channel ==6'b000000) nextState=ch0;
else if (channel ==6'b011100) nextState=ch28;
else if (channel ==6'b011101) nextState=ch29;
else if (channel ==6'b011110) nextState=ch30;
else if (channel ==6'b011111) nextState=ch31;
else if (channel ==6'b100000) nextState=ch32;
else if (channel ==6'b100001) nextState=ch33;
else if (channel ==6'b100010) nextState=ch34;
else if (channel ==6'b100011) nextState=ch35;
else if (channel ==6'b100100) nextState=ch36;
else if (channel ==6'b100101) nextState=ch37;
else if (channel ==6'b100110) nextState=ch38;
else if (channel ==6'b100111) nextState=ch39;
else if (channel ==6'b101000) nextState=ch40;
else if (channel ==6'b101001) nextState=ch41;
else if (channel ==6'b101010) nextState=ch42;
else if (channel ==6'b101011) nextState=ch43;
else if (channel ==6'b101100) nextState=ch44;
else if (channel ==6'b101101) nextState=ch45;
else if (channel ==6'b101110) nextState=ch46;
else if (channel ==6'b101111) nextState=ch47;
else if (channel ==6'b110000) nextState=ch48;
else if (channel ==6'b110001) nextState=ch49;
else if (channel ==6'b110010) nextState=ch50;
else if (channel ==6'b110011) nextState=ch51;
else if (channel ==6'b110100) nextState=ch52;
else if (channel ==6'b110101) nextState=ch53;
else if (channel ==6'b110110) nextState=ch54;
else if (channel ==6'b110111) nextState=ch55;
else if (channel ==6'b111000) nextState=ch56;
else if (channel ==6'b111001) nextState=ch57;
else if (channel ==6'b111010) nextState=ch58;
else if (channel ==6'b111011) nextState=ch59;
else if (channel ==6'b111100) nextState=ch60;
else if (channel ==6'b111101) nextState=ch61;
else if (channel ==6'b111110) nextState=ch62;
else nextState=ch63;


ch28:if (channel ==6'b011100) nextState=ch28;
else if (channel ==6'b000001) nextState=ch1;
else if (channel ==6'b000010) nextState=ch2;
else if (channel ==6'b000011) nextState=ch3;
else if (channel ==6'b000100) nextState=ch4;
else if (channel ==6'b000101) nextState=ch5;
else if (channel ==6'b000110) nextState=ch6;
else if (channel ==6'b000111) nextState=ch7;
else if (channel ==6'b001000) nextState=ch8;
else if (channel ==6'b001001) nextState=ch9;
else if (channel ==6'b001010) nextState=ch10;
else if (channel ==6'b001011) nextState=ch11;
else if (channel ==6'b001100) nextState=ch12;
else if (channel ==6'b001101) nextState=ch13;
else if (channel ==6'b001110) nextState=ch14;
else if (channel ==6'b001111) nextState=ch15;
else if (channel ==6'b010000) nextState=ch16;
else if (channel ==6'b010001) nextState=ch17;
else if (channel ==6'b010010) nextState=ch18;
else if (channel ==6'b010011) nextState=ch19;
else if (channel ==6'b010100) nextState=ch20;
else if (channel ==6'b010101) nextState=ch21;
else if (channel ==6'b010110) nextState=ch22;
else if (channel ==6'b010111) nextState=ch23;
else if (channel ==6'b011000) nextState=ch24;
else if (channel ==6'b011001) nextState=ch25;
else if (channel ==6'b011010) nextState=ch26;
else if (channel ==6'b011011) nextState=ch27;
else if (channel ==6'b000000) nextState=ch0;
else if (channel ==6'b011101) nextState=ch29;
else if (channel ==6'b011110) nextState=ch30;
else if (channel ==6'b011111) nextState=ch31;
else if (channel ==6'b100000) nextState=ch32;
else if (channel ==6'b100001) nextState=ch33;
else if (channel ==6'b100010) nextState=ch34;
else if (channel ==6'b100011) nextState=ch35;
else if (channel ==6'b100100) nextState=ch36;
else if (channel ==6'b100101) nextState=ch37;
else if (channel ==6'b100110) nextState=ch38;
else if (channel ==6'b100111) nextState=ch39;
else if (channel ==6'b101000) nextState=ch40;
else if (channel ==6'b101001) nextState=ch41;
else if (channel ==6'b101010) nextState=ch42;
else if (channel ==6'b101011) nextState=ch43;
else if (channel ==6'b101100) nextState=ch44;
else if (channel ==6'b101101) nextState=ch45;
else if (channel ==6'b101110) nextState=ch46;
else if (channel ==6'b101111) nextState=ch47;
else if (channel ==6'b110000) nextState=ch48;
else if (channel ==6'b110001) nextState=ch49;
else if (channel ==6'b110010) nextState=ch50;
else if (channel ==6'b110011) nextState=ch51;
else if (channel ==6'b110100) nextState=ch52;
else if (channel ==6'b110101) nextState=ch53;
else if (channel ==6'b110110) nextState=ch54;
else if (channel ==6'b110111) nextState=ch55;
else if (channel ==6'b111000) nextState=ch56;
else if (channel ==6'b111001) nextState=ch57;
else if (channel ==6'b111010) nextState=ch58;
else if (channel ==6'b111011) nextState=ch59;
else if (channel ==6'b111100) nextState=ch60;
else if (channel ==6'b111101) nextState=ch61;
else if (channel ==6'b111110) nextState=ch62;
else nextState=ch63;


ch29:if (channel ==6'b011101) nextState=ch29;
else if (channel ==6'b000001) nextState=ch1;
else if (channel ==6'b000010) nextState=ch2;
else if (channel ==6'b000011) nextState=ch3;
else if (channel ==6'b000100) nextState=ch4;
else if (channel ==6'b000101) nextState=ch5;
else if (channel ==6'b000110) nextState=ch6;
else if (channel ==6'b000111) nextState=ch7;
else if (channel ==6'b001000) nextState=ch8;
else if (channel ==6'b001001) nextState=ch9;
else if (channel ==6'b001010) nextState=ch10;
else if (channel ==6'b001011) nextState=ch11;
else if (channel ==6'b001100) nextState=ch12;
else if (channel ==6'b001101) nextState=ch13;
else if (channel ==6'b001110) nextState=ch14;
else if (channel ==6'b001111) nextState=ch15;
else if (channel ==6'b010000) nextState=ch16;
else if (channel ==6'b010001) nextState=ch17;
else if (channel ==6'b010010) nextState=ch18;
else if (channel ==6'b010011) nextState=ch19;
else if (channel ==6'b010100) nextState=ch20;
else if (channel ==6'b010101) nextState=ch21;
else if (channel ==6'b010110) nextState=ch22;
else if (channel ==6'b010111) nextState=ch23;
else if (channel ==6'b011000) nextState=ch24;
else if (channel ==6'b011001) nextState=ch25;
else if (channel ==6'b011010) nextState=ch26;
else if (channel ==6'b011011) nextState=ch27;
else if (channel ==6'b011100) nextState=ch28;
else if (channel ==6'b000000) nextState=ch0;
else if (channel ==6'b011110) nextState=ch30;
else if (channel ==6'b011111) nextState=ch31;
else if (channel ==6'b100000) nextState=ch32;
else if (channel ==6'b100001) nextState=ch33;
else if (channel ==6'b100010) nextState=ch34;
else if (channel ==6'b100011) nextState=ch35;
else if (channel ==6'b100100) nextState=ch36;
else if (channel ==6'b100101) nextState=ch37;
else if (channel ==6'b100110) nextState=ch38;
else if (channel ==6'b100111) nextState=ch39;
else if (channel ==6'b101000) nextState=ch40;
else if (channel ==6'b101001) nextState=ch41;
else if (channel ==6'b101010) nextState=ch42;
else if (channel ==6'b101011) nextState=ch43;
else if (channel ==6'b101100) nextState=ch44;
else if (channel ==6'b101101) nextState=ch45;
else if (channel ==6'b101110) nextState=ch46;
else if (channel ==6'b101111) nextState=ch47;
else if (channel ==6'b110000) nextState=ch48;
else if (channel ==6'b110001) nextState=ch49;
else if (channel ==6'b110010) nextState=ch50;
else if (channel ==6'b110011) nextState=ch51;
else if (channel ==6'b110100) nextState=ch52;
else if (channel ==6'b110101) nextState=ch53;
else if (channel ==6'b110110) nextState=ch54;
else if (channel ==6'b110111) nextState=ch55;
else if (channel ==6'b111000) nextState=ch56;
else if (channel ==6'b111001) nextState=ch57;
else if (channel ==6'b111010) nextState=ch58;
else if (channel ==6'b111011) nextState=ch59;
else if (channel ==6'b111100) nextState=ch60;
else if (channel ==6'b111101) nextState=ch61;
else if (channel ==6'b111110) nextState=ch62;
else nextState=ch63;


ch30:if (channel ==6'b011110) nextState=ch30;
else if (channel ==6'b000001) nextState=ch1;
else if (channel ==6'b000010) nextState=ch2;
else if (channel ==6'b000011) nextState=ch3;
else if (channel ==6'b000100) nextState=ch4;
else if (channel ==6'b000101) nextState=ch5;
else if (channel ==6'b000110) nextState=ch6;
else if (channel ==6'b000111) nextState=ch7;
else if (channel ==6'b001000) nextState=ch8;
else if (channel ==6'b001001) nextState=ch9;
else if (channel ==6'b001010) nextState=ch10;
else if (channel ==6'b001011) nextState=ch11;
else if (channel ==6'b001100) nextState=ch12;
else if (channel ==6'b001101) nextState=ch13;
else if (channel ==6'b001110) nextState=ch14;
else if (channel ==6'b001111) nextState=ch15;
else if (channel ==6'b010000) nextState=ch16;
else if (channel ==6'b010001) nextState=ch17;
else if (channel ==6'b010010) nextState=ch18;
else if (channel ==6'b010011) nextState=ch19;
else if (channel ==6'b010100) nextState=ch20;
else if (channel ==6'b010101) nextState=ch21;
else if (channel ==6'b010110) nextState=ch22;
else if (channel ==6'b010111) nextState=ch23;
else if (channel ==6'b011000) nextState=ch24;
else if (channel ==6'b011001) nextState=ch25;
else if (channel ==6'b011010) nextState=ch26;
else if (channel ==6'b011011) nextState=ch27;
else if (channel ==6'b011100) nextState=ch28;
else if (channel ==6'b011101) nextState=ch29;
else if (channel ==6'b000000) nextState=ch0;
else if (channel ==6'b011111) nextState=ch31;
else if (channel ==6'b100000) nextState=ch32;
else if (channel ==6'b100001) nextState=ch33;
else if (channel ==6'b100010) nextState=ch34;
else if (channel ==6'b100011) nextState=ch35;
else if (channel ==6'b100100) nextState=ch36;
else if (channel ==6'b100101) nextState=ch37;
else if (channel ==6'b100110) nextState=ch38;
else if (channel ==6'b100111) nextState=ch39;
else if (channel ==6'b101000) nextState=ch40;
else if (channel ==6'b101001) nextState=ch41;
else if (channel ==6'b101010) nextState=ch42;
else if (channel ==6'b101011) nextState=ch43;
else if (channel ==6'b101100) nextState=ch44;
else if (channel ==6'b101101) nextState=ch45;
else if (channel ==6'b101110) nextState=ch46;
else if (channel ==6'b101111) nextState=ch47;
else if (channel ==6'b110000) nextState=ch48;
else if (channel ==6'b110001) nextState=ch49;
else if (channel ==6'b110010) nextState=ch50;
else if (channel ==6'b110011) nextState=ch51;
else if (channel ==6'b110100) nextState=ch52;
else if (channel ==6'b110101) nextState=ch53;
else if (channel ==6'b110110) nextState=ch54;
else if (channel ==6'b110111) nextState=ch55;
else if (channel ==6'b111000) nextState=ch56;
else if (channel ==6'b111001) nextState=ch57;
else if (channel ==6'b111010) nextState=ch58;
else if (channel ==6'b111011) nextState=ch59;
else if (channel ==6'b111100) nextState=ch60;
else if (channel ==6'b111101) nextState=ch61;
else if (channel ==6'b111110) nextState=ch62;
else nextState=ch63;


ch31:if (channel ==5'b11111) nextState=ch31;
else if (channel ==6'b000001) nextState=ch1;
else if (channel ==6'b000010) nextState=ch2;
else if (channel ==6'b000011) nextState=ch3;
else if (channel ==6'b000100) nextState=ch4;
else if (channel ==6'b000101) nextState=ch5;
else if (channel ==6'b000110) nextState=ch6;
else if (channel ==6'b000111) nextState=ch7;
else if (channel ==6'b001000) nextState=ch8;
else if (channel ==6'b001001) nextState=ch9;
else if (channel ==6'b001010) nextState=ch10;
else if (channel ==6'b001011) nextState=ch11;
else if (channel ==6'b001100) nextState=ch12;
else if (channel ==6'b001101) nextState=ch13;
else if (channel ==6'b001110) nextState=ch14;
else if (channel ==6'b001111) nextState=ch15;
else if (channel ==6'b010000) nextState=ch16;
else if (channel ==6'b010001) nextState=ch17;
else if (channel ==6'b010010) nextState=ch18;
else if (channel ==6'b010011) nextState=ch19;
else if (channel ==6'b010100) nextState=ch20;
else if (channel ==6'b010101) nextState=ch21;
else if (channel ==6'b010110) nextState=ch22;
else if (channel ==6'b010111) nextState=ch23;
else if (channel ==6'b011000) nextState=ch24;
else if (channel ==6'b011001) nextState=ch25;
else if (channel ==6'b011010) nextState=ch26;
else if (channel ==6'b011011) nextState=ch27;
else if (channel ==6'b011100) nextState=ch28;
else if (channel ==6'b011101) nextState=ch29;
else if (channel ==6'b011110) nextState=ch30;
else if (channel == 6'b000000) nextState=ch0;
else if (channel ==6'b100000) nextState=ch32;
else if (channel ==6'b100001) nextState=ch33;
else if (channel ==6'b100010) nextState=ch34;
else if (channel ==6'b100011) nextState=ch35;
else if (channel ==6'b100100) nextState=ch36;
else if (channel ==6'b100101) nextState=ch37;
else if (channel ==6'b100110) nextState=ch38;
else if (channel ==6'b100111) nextState=ch39;
else if (channel ==6'b101000) nextState=ch40;
else if (channel ==6'b101001) nextState=ch41;
else if (channel ==6'b101010) nextState=ch42;
else if (channel ==6'b101011) nextState=ch43;
else if (channel ==6'b101100) nextState=ch44;
else if (channel ==6'b101101) nextState=ch45;
else if (channel ==6'b101110) nextState=ch46;
else if (channel ==6'b101111) nextState=ch47;
else if (channel ==6'b110000) nextState=ch48;
else if (channel ==6'b110001) nextState=ch49;
else if (channel ==6'b110010) nextState=ch50;
else if (channel ==6'b110011) nextState=ch51;
else if (channel ==6'b110100) nextState=ch52;
else if (channel ==6'b110101) nextState=ch53;
else if (channel ==6'b110110) nextState=ch54;
else if (channel ==6'b110111) nextState=ch55;
else if (channel ==6'b111000) nextState=ch56;
else if (channel ==6'b111001) nextState=ch57;
else if (channel ==6'b111010) nextState=ch58;
else if (channel ==6'b111011) nextState=ch59;
else if (channel ==6'b111100) nextState=ch60;
else if (channel ==6'b111101) nextState=ch61;
else if (channel ==6'b111110) nextState=ch62;
else nextState=ch63;

ch32: 
if (channel == 6'b100000) nextState=ch32;
else if (channel ==6'b000001) nextState=ch1;
else if (channel ==6'b000010) nextState=ch2;
else if (channel ==6'b000011) nextState=ch3;
else if (channel ==6'b000100) nextState=ch4;
else if (channel ==6'b000101) nextState=ch5;
else if (channel ==6'b000110) nextState=ch6;
else if (channel ==6'b000111) nextState=ch7;
else if (channel ==6'b001000) nextState=ch8;
else if (channel ==6'b001001) nextState=ch9;
else if (channel ==6'b001010) nextState=ch10;
else if (channel ==6'b001011) nextState=ch11;
else if (channel ==6'b001100) nextState=ch12;
else if (channel ==6'b001101) nextState=ch13;
else if (channel ==6'b001110) nextState=ch14;
else if (channel ==6'b001111) nextState=ch15;
else if (channel ==6'b010000) nextState=ch16;
else if (channel ==6'b010001) nextState=ch17;
else if (channel ==6'b010010) nextState=ch18;
else if (channel ==6'b010011) nextState=ch19;
else if (channel ==6'b010100) nextState=ch20;
else if (channel ==6'b010101) nextState=ch21;
else if (channel ==6'b010110) nextState=ch22;
else if (channel ==6'b010111) nextState=ch23;
else if (channel ==6'b011000) nextState=ch24;
else if (channel ==6'b011001) nextState=ch25;
else if (channel ==6'b011010) nextState=ch26;
else if (channel ==6'b011011) nextState=ch27;
else if (channel ==6'b011100) nextState=ch28;
else if (channel ==6'b011101) nextState=ch29;
else if (channel ==6'b011110) nextState=ch30;
else if (channel ==6'b011111) nextState=ch31;
else if (channel ==6'b000000) nextState=ch0;
else if (channel ==6'b100001) nextState=ch33;
else if (channel ==6'b100010) nextState=ch34;
else if (channel ==6'b100011) nextState=ch35;
else if (channel ==6'b100100) nextState=ch36;
else if (channel ==6'b100101) nextState=ch37;
else if (channel ==6'b100110) nextState=ch38;
else if (channel ==6'b100111) nextState=ch39;
else if (channel ==6'b101000) nextState=ch40;
else if (channel ==6'b101001) nextState=ch41;
else if (channel ==6'b101010) nextState=ch42;
else if (channel ==6'b101011) nextState=ch43;
else if (channel ==6'b101100) nextState=ch44;
else if (channel ==6'b101101) nextState=ch45;
else if (channel ==6'b101110) nextState=ch46;
else if (channel ==6'b101111) nextState=ch47;
else if (channel ==6'b110000) nextState=ch48;
else if (channel ==6'b110001) nextState=ch49;
else if (channel ==6'b110010) nextState=ch50;
else if (channel ==6'b110011) nextState=ch51;
else if (channel ==6'b110100) nextState=ch52;
else if (channel ==6'b110101) nextState=ch53;
else if (channel ==6'b110110) nextState=ch54;
else if (channel ==6'b110111) nextState=ch55;
else if (channel ==6'b111000) nextState=ch56;
else if (channel ==6'b111001) nextState=ch57;
else if (channel ==6'b111010) nextState=ch58;
else if (channel ==6'b111011) nextState=ch59;
else if (channel ==6'b111100) nextState=ch60;
else if (channel ==6'b111101) nextState=ch61;
else if (channel ==6'b111110) nextState=ch62;
else nextState=ch63;

ch33: 
if (channel == 6'b100001) nextState=ch33;
else if (channel ==6'b000001) nextState=ch1;
else if (channel ==6'b000010) nextState=ch2;
else if (channel ==6'b000011) nextState=ch3;
else if (channel ==6'b000100) nextState=ch4;
else if (channel ==6'b000101) nextState=ch5;
else if (channel ==6'b000110) nextState=ch6;
else if (channel ==6'b000111) nextState=ch7;
else if (channel ==6'b001000) nextState=ch8;
else if (channel ==6'b001001) nextState=ch9;
else if (channel ==6'b001010) nextState=ch10;
else if (channel ==6'b001011) nextState=ch11;
else if (channel ==6'b001100) nextState=ch12;
else if (channel ==6'b001101) nextState=ch13;
else if (channel ==6'b001110) nextState=ch14;
else if (channel ==6'b001111) nextState=ch15;
else if (channel ==6'b010000) nextState=ch16;
else if (channel ==6'b010001) nextState=ch17;
else if (channel ==6'b010010) nextState=ch18;
else if (channel ==6'b010011) nextState=ch19;
else if (channel ==6'b010100) nextState=ch20;
else if (channel ==6'b010101) nextState=ch21;
else if (channel ==6'b010110) nextState=ch22;
else if (channel ==6'b010111) nextState=ch23;
else if (channel ==6'b011000) nextState=ch24;
else if (channel ==6'b011001) nextState=ch25;
else if (channel ==6'b011010) nextState=ch26;
else if (channel ==6'b011011) nextState=ch27;
else if (channel ==6'b011100) nextState=ch28;
else if (channel ==6'b011101) nextState=ch29;
else if (channel ==6'b011110) nextState=ch30;
else if (channel ==6'b011111) nextState=ch31;
else if (channel ==6'b100000) nextState=ch32;
else if (channel ==6'b000000) nextState=ch0;
else if (channel ==6'b100010) nextState=ch34;
else if (channel ==6'b100011) nextState=ch35;
else if (channel ==6'b100100) nextState=ch36;
else if (channel ==6'b100101) nextState=ch37;
else if (channel ==6'b100110) nextState=ch38;
else if (channel ==6'b100111) nextState=ch39;
else if (channel ==6'b101000) nextState=ch40;
else if (channel ==6'b101001) nextState=ch41;
else if (channel ==6'b101010) nextState=ch42;
else if (channel ==6'b101011) nextState=ch43;
else if (channel ==6'b101100) nextState=ch44;
else if (channel ==6'b101101) nextState=ch45;
else if (channel ==6'b101110) nextState=ch46;
else if (channel ==6'b101111) nextState=ch47;
else if (channel ==6'b110000) nextState=ch48;
else if (channel ==6'b110001) nextState=ch49;
else if (channel ==6'b110010) nextState=ch50;
else if (channel ==6'b110011) nextState=ch51;
else if (channel ==6'b110100) nextState=ch52;
else if (channel ==6'b110101) nextState=ch53;
else if (channel ==6'b110110) nextState=ch54;
else if (channel ==6'b110111) nextState=ch55;
else if (channel ==6'b111000) nextState=ch56;
else if (channel ==6'b111001) nextState=ch57;
else if (channel ==6'b111010) nextState=ch58;
else if (channel ==6'b111011) nextState=ch59;
else if (channel ==6'b111100) nextState=ch60;
else if (channel ==6'b111101) nextState=ch61;
else if (channel ==6'b111110) nextState=ch62;
else nextState=ch63;

ch34: 
if (channel == 6'b100010) nextState=ch34;
else if (channel ==6'b000001) nextState=ch1;
else if (channel ==6'b000010) nextState=ch2;
else if (channel ==6'b000011) nextState=ch3;
else if (channel ==6'b000100) nextState=ch4;
else if (channel ==6'b000101) nextState=ch5;
else if (channel ==6'b000110) nextState=ch6;
else if (channel ==6'b000111) nextState=ch7;
else if (channel ==6'b001000) nextState=ch8;
else if (channel ==6'b001001) nextState=ch9;
else if (channel ==6'b001010) nextState=ch10;
else if (channel ==6'b001011) nextState=ch11;
else if (channel ==6'b001100) nextState=ch12;
else if (channel ==6'b001101) nextState=ch13;
else if (channel ==6'b001110) nextState=ch14;
else if (channel ==6'b001111) nextState=ch15;
else if (channel ==6'b010000) nextState=ch16;
else if (channel ==6'b010001) nextState=ch17;
else if (channel ==6'b010010) nextState=ch18;
else if (channel ==6'b010011) nextState=ch19;
else if (channel ==6'b010100) nextState=ch20;
else if (channel ==6'b010101) nextState=ch21;
else if (channel ==6'b010110) nextState=ch22;
else if (channel ==6'b010111) nextState=ch23;
else if (channel ==6'b011000) nextState=ch24;
else if (channel ==6'b011001) nextState=ch25;
else if (channel ==6'b011010) nextState=ch26;
else if (channel ==6'b011011) nextState=ch27;
else if (channel ==6'b011100) nextState=ch28;
else if (channel ==6'b011101) nextState=ch29;
else if (channel ==6'b011110) nextState=ch30;
else if (channel ==6'b011111) nextState=ch31;
else if (channel ==6'b100000) nextState=ch32;
else if (channel ==6'b100001) nextState=ch33;
else if (channel ==6'b000000) nextState=ch0;
else if (channel ==6'b100011) nextState=ch35;
else if (channel ==6'b100100) nextState=ch36;
else if (channel ==6'b100101) nextState=ch37;
else if (channel ==6'b100110) nextState=ch38;
else if (channel ==6'b100111) nextState=ch39;
else if (channel ==6'b101000) nextState=ch40;
else if (channel ==6'b101001) nextState=ch41;
else if (channel ==6'b101010) nextState=ch42;
else if (channel ==6'b101011) nextState=ch43;
else if (channel ==6'b101100) nextState=ch44;
else if (channel ==6'b101101) nextState=ch45;
else if (channel ==6'b101110) nextState=ch46;
else if (channel ==6'b101111) nextState=ch47;
else if (channel ==6'b110000) nextState=ch48;
else if (channel ==6'b110001) nextState=ch49;
else if (channel ==6'b110010) nextState=ch50;
else if (channel ==6'b110011) nextState=ch51;
else if (channel ==6'b110100) nextState=ch52;
else if (channel ==6'b110101) nextState=ch53;
else if (channel ==6'b110110) nextState=ch54;
else if (channel ==6'b110111) nextState=ch55;
else if (channel ==6'b111000) nextState=ch56;
else if (channel ==6'b111001) nextState=ch57;
else if (channel ==6'b111010) nextState=ch58;
else if (channel ==6'b111011) nextState=ch59;
else if (channel ==6'b111100) nextState=ch60;
else if (channel ==6'b111101) nextState=ch61;
else if (channel ==6'b111110) nextState=ch62;
else nextState=ch63;

ch35: 
if (channel == 6'b100011) nextState=ch35;
else if (channel ==6'b000001) nextState=ch1;
else if (channel ==6'b000010) nextState=ch2;
else if (channel ==6'b000011) nextState=ch3;
else if (channel ==6'b000100) nextState=ch4;
else if (channel ==6'b000101) nextState=ch5;
else if (channel ==6'b000110) nextState=ch6;
else if (channel ==6'b000111) nextState=ch7;
else if (channel ==6'b001000) nextState=ch8;
else if (channel ==6'b001001) nextState=ch9;
else if (channel ==6'b001010) nextState=ch10;
else if (channel ==6'b001011) nextState=ch11;
else if (channel ==6'b001100) nextState=ch12;
else if (channel ==6'b001101) nextState=ch13;
else if (channel ==6'b001110) nextState=ch14;
else if (channel ==6'b001111) nextState=ch15;
else if (channel ==6'b010000) nextState=ch16;
else if (channel ==6'b010001) nextState=ch17;
else if (channel ==6'b010010) nextState=ch18;
else if (channel ==6'b010011) nextState=ch19;
else if (channel ==6'b010100) nextState=ch20;
else if (channel ==6'b010101) nextState=ch21;
else if (channel ==6'b010110) nextState=ch22;
else if (channel ==6'b010111) nextState=ch23;
else if (channel ==6'b011000) nextState=ch24;
else if (channel ==6'b011001) nextState=ch25;
else if (channel ==6'b011010) nextState=ch26;
else if (channel ==6'b011011) nextState=ch27;
else if (channel ==6'b011100) nextState=ch28;
else if (channel ==6'b011101) nextState=ch29;
else if (channel ==6'b011110) nextState=ch30;
else if (channel ==6'b011111) nextState=ch31;
else if (channel ==6'b100000) nextState=ch32;
else if (channel ==6'b100001) nextState=ch33;
else if (channel ==6'b100010) nextState=ch34;
else if (channel ==6'b000000) nextState=ch0;
else if (channel ==6'b100100) nextState=ch36;
else if (channel ==6'b100101) nextState=ch37;
else if (channel ==6'b100110) nextState=ch38;
else if (channel ==6'b100111) nextState=ch39;
else if (channel ==6'b101000) nextState=ch40;
else if (channel ==6'b101001) nextState=ch41;
else if (channel ==6'b101010) nextState=ch42;
else if (channel ==6'b101011) nextState=ch43;
else if (channel ==6'b101100) nextState=ch44;
else if (channel ==6'b101101) nextState=ch45;
else if (channel ==6'b101110) nextState=ch46;
else if (channel ==6'b101111) nextState=ch47;
else if (channel ==6'b110000) nextState=ch48;
else if (channel ==6'b110001) nextState=ch49;
else if (channel ==6'b110010) nextState=ch50;
else if (channel ==6'b110011) nextState=ch51;
else if (channel ==6'b110100) nextState=ch52;
else if (channel ==6'b110101) nextState=ch53;
else if (channel ==6'b110110) nextState=ch54;
else if (channel ==6'b110111) nextState=ch55;
else if (channel ==6'b111000) nextState=ch56;
else if (channel ==6'b111001) nextState=ch57;
else if (channel ==6'b111010) nextState=ch58;
else if (channel ==6'b111011) nextState=ch59;
else if (channel ==6'b111100) nextState=ch60;
else if (channel ==6'b111101) nextState=ch61;
else if (channel ==6'b111110) nextState=ch62;
else nextState=ch63;

ch36: 
if (channel == 6'b100100) nextState=ch36;
else if (channel ==6'b000001) nextState=ch1;
else if (channel ==6'b000010) nextState=ch2;
else if (channel ==6'b000011) nextState=ch3;
else if (channel ==6'b000100) nextState=ch4;
else if (channel ==6'b000101) nextState=ch5;
else if (channel ==6'b000110) nextState=ch6;
else if (channel ==6'b000111) nextState=ch7;
else if (channel ==6'b001000) nextState=ch8;
else if (channel ==6'b001001) nextState=ch9;
else if (channel ==6'b001010) nextState=ch10;
else if (channel ==6'b001011) nextState=ch11;
else if (channel ==6'b001100) nextState=ch12;
else if (channel ==6'b001101) nextState=ch13;
else if (channel ==6'b001110) nextState=ch14;
else if (channel ==6'b001111) nextState=ch15;
else if (channel ==6'b010000) nextState=ch16;
else if (channel ==6'b010001) nextState=ch17;
else if (channel ==6'b010010) nextState=ch18;
else if (channel ==6'b010011) nextState=ch19;
else if (channel ==6'b010100) nextState=ch20;
else if (channel ==6'b010101) nextState=ch21;
else if (channel ==6'b010110) nextState=ch22;
else if (channel ==6'b010111) nextState=ch23;
else if (channel ==6'b011000) nextState=ch24;
else if (channel ==6'b011001) nextState=ch25;
else if (channel ==6'b011010) nextState=ch26;
else if (channel ==6'b011011) nextState=ch27;
else if (channel ==6'b011100) nextState=ch28;
else if (channel ==6'b011101) nextState=ch29;
else if (channel ==6'b011110) nextState=ch30;
else if (channel ==6'b011111) nextState=ch31;
else if (channel ==6'b100000) nextState=ch32;
else if (channel ==6'b100001) nextState=ch33;
else if (channel ==6'b100010) nextState=ch34;
else if (channel ==6'b100011) nextState=ch35;
else if (channel ==6'b000000) nextState=ch0;
else if (channel ==6'b100101) nextState=ch37;
else if (channel ==6'b100110) nextState=ch38;
else if (channel ==6'b100111) nextState=ch39;
else if (channel ==6'b101000) nextState=ch40;
else if (channel ==6'b101001) nextState=ch41;
else if (channel ==6'b101010) nextState=ch42;
else if (channel ==6'b101011) nextState=ch43;
else if (channel ==6'b101100) nextState=ch44;
else if (channel ==6'b101101) nextState=ch45;
else if (channel ==6'b101110) nextState=ch46;
else if (channel ==6'b101111) nextState=ch47;
else if (channel ==6'b110000) nextState=ch48;
else if (channel ==6'b110001) nextState=ch49;
else if (channel ==6'b110010) nextState=ch50;
else if (channel ==6'b110011) nextState=ch51;
else if (channel ==6'b110100) nextState=ch52;
else if (channel ==6'b110101) nextState=ch53;
else if (channel ==6'b110110) nextState=ch54;
else if (channel ==6'b110111) nextState=ch55;
else if (channel ==6'b111000) nextState=ch56;
else if (channel ==6'b111001) nextState=ch57;
else if (channel ==6'b111010) nextState=ch58;
else if (channel ==6'b111011) nextState=ch59;
else if (channel ==6'b111100) nextState=ch60;
else if (channel ==6'b111101) nextState=ch61;
else if (channel ==6'b111110) nextState=ch62;
else nextState=ch63;

ch37: 
if (channel == 6'b100101) nextState=ch37;
else if (channel ==6'b000001) nextState=ch1;
else if (channel ==6'b000010) nextState=ch2;
else if (channel ==6'b000011) nextState=ch3;
else if (channel ==6'b000100) nextState=ch4;
else if (channel ==6'b000101) nextState=ch5;
else if (channel ==6'b000110) nextState=ch6;
else if (channel ==6'b000111) nextState=ch7;
else if (channel ==6'b001000) nextState=ch8;
else if (channel ==6'b001001) nextState=ch9;
else if (channel ==6'b001010) nextState=ch10;
else if (channel ==6'b001011) nextState=ch11;
else if (channel ==6'b001100) nextState=ch12;
else if (channel ==6'b001101) nextState=ch13;
else if (channel ==6'b001110) nextState=ch14;
else if (channel ==6'b001111) nextState=ch15;
else if (channel ==6'b010000) nextState=ch16;
else if (channel ==6'b010001) nextState=ch17;
else if (channel ==6'b010010) nextState=ch18;
else if (channel ==6'b010011) nextState=ch19;
else if (channel ==6'b010100) nextState=ch20;
else if (channel ==6'b010101) nextState=ch21;
else if (channel ==6'b010110) nextState=ch22;
else if (channel ==6'b010111) nextState=ch23;
else if (channel ==6'b011000) nextState=ch24;
else if (channel ==6'b011001) nextState=ch25;
else if (channel ==6'b011010) nextState=ch26;
else if (channel ==6'b011011) nextState=ch27;
else if (channel ==6'b011100) nextState=ch28;
else if (channel ==6'b011101) nextState=ch29;
else if (channel ==6'b011110) nextState=ch30;
else if (channel ==6'b011111) nextState=ch31;
else if (channel ==6'b100000) nextState=ch32;
else if (channel ==6'b100001) nextState=ch33;
else if (channel ==6'b100010) nextState=ch34;
else if (channel ==6'b100011) nextState=ch35;
else if (channel ==6'b100100) nextState=ch36;
else if (channel ==6'b000000) nextState=ch0;
else if (channel ==6'b100110) nextState=ch38;
else if (channel ==6'b100111) nextState=ch39;
else if (channel ==6'b101000) nextState=ch40;
else if (channel ==6'b101001) nextState=ch41;
else if (channel ==6'b101010) nextState=ch42;
else if (channel ==6'b101011) nextState=ch43;
else if (channel ==6'b101100) nextState=ch44;
else if (channel ==6'b101101) nextState=ch45;
else if (channel ==6'b101110) nextState=ch46;
else if (channel ==6'b101111) nextState=ch47;
else if (channel ==6'b110000) nextState=ch48;
else if (channel ==6'b110001) nextState=ch49;
else if (channel ==6'b110010) nextState=ch50;
else if (channel ==6'b110011) nextState=ch51;
else if (channel ==6'b110100) nextState=ch52;
else if (channel ==6'b110101) nextState=ch53;
else if (channel ==6'b110110) nextState=ch54;
else if (channel ==6'b110111) nextState=ch55;
else if (channel ==6'b111000) nextState=ch56;
else if (channel ==6'b111001) nextState=ch57;
else if (channel ==6'b111010) nextState=ch58;
else if (channel ==6'b111011) nextState=ch59;
else if (channel ==6'b111100) nextState=ch60;
else if (channel ==6'b111101) nextState=ch61;
else if (channel ==6'b111110) nextState=ch62;
else nextState=ch63;

ch38: 
if (channel == 6'b100110) nextState=ch38;
else if (channel ==6'b000001) nextState=ch1;
else if (channel ==6'b000010) nextState=ch2;
else if (channel ==6'b000011) nextState=ch3;
else if (channel ==6'b000100) nextState=ch4;
else if (channel ==6'b000101) nextState=ch5;
else if (channel ==6'b000110) nextState=ch6;
else if (channel ==6'b000111) nextState=ch7;
else if (channel ==6'b001000) nextState=ch8;
else if (channel ==6'b001001) nextState=ch9;
else if (channel ==6'b001010) nextState=ch10;
else if (channel ==6'b001011) nextState=ch11;
else if (channel ==6'b001100) nextState=ch12;
else if (channel ==6'b001101) nextState=ch13;
else if (channel ==6'b001110) nextState=ch14;
else if (channel ==6'b001111) nextState=ch15;
else if (channel ==6'b010000) nextState=ch16;
else if (channel ==6'b010001) nextState=ch17;
else if (channel ==6'b010010) nextState=ch18;
else if (channel ==6'b010011) nextState=ch19;
else if (channel ==6'b010100) nextState=ch20;
else if (channel ==6'b010101) nextState=ch21;
else if (channel ==6'b010110) nextState=ch22;
else if (channel ==6'b010111) nextState=ch23;
else if (channel ==6'b011000) nextState=ch24;
else if (channel ==6'b011001) nextState=ch25;
else if (channel ==6'b011010) nextState=ch26;
else if (channel ==6'b011011) nextState=ch27;
else if (channel ==6'b011100) nextState=ch28;
else if (channel ==6'b011101) nextState=ch29;
else if (channel ==6'b011110) nextState=ch30;
else if (channel ==6'b011111) nextState=ch31;
else if (channel ==6'b100000) nextState=ch32;
else if (channel ==6'b100001) nextState=ch33;
else if (channel ==6'b100010) nextState=ch34;
else if (channel ==6'b100011) nextState=ch35;
else if (channel ==6'b100100) nextState=ch36;
else if (channel ==6'b100101) nextState=ch37;
else if (channel ==6'b000000) nextState=ch0;
else if (channel ==6'b100111) nextState=ch39;
else if (channel ==6'b101000) nextState=ch40;
else if (channel ==6'b101001) nextState=ch41;
else if (channel ==6'b101010) nextState=ch42;
else if (channel ==6'b101011) nextState=ch43;
else if (channel ==6'b101100) nextState=ch44;
else if (channel ==6'b101101) nextState=ch45;
else if (channel ==6'b101110) nextState=ch46;
else if (channel ==6'b101111) nextState=ch47;
else if (channel ==6'b110000) nextState=ch48;
else if (channel ==6'b110001) nextState=ch49;
else if (channel ==6'b110010) nextState=ch50;
else if (channel ==6'b110011) nextState=ch51;
else if (channel ==6'b110100) nextState=ch52;
else if (channel ==6'b110101) nextState=ch53;
else if (channel ==6'b110110) nextState=ch54;
else if (channel ==6'b110111) nextState=ch55;
else if (channel ==6'b111000) nextState=ch56;
else if (channel ==6'b111001) nextState=ch57;
else if (channel ==6'b111010) nextState=ch58;
else if (channel ==6'b111011) nextState=ch59;
else if (channel ==6'b111100) nextState=ch60;
else if (channel ==6'b111101) nextState=ch61;
else if (channel ==6'b111110) nextState=ch62;
else nextState=ch63;

ch39: 
if (channel == 6'b100111) nextState=ch39;
else if (channel ==6'b000001) nextState=ch1;
else if (channel ==6'b000010) nextState=ch2;
else if (channel ==6'b000011) nextState=ch3;
else if (channel ==6'b000100) nextState=ch4;
else if (channel ==6'b000101) nextState=ch5;
else if (channel ==6'b000110) nextState=ch6;
else if (channel ==6'b000111) nextState=ch7;
else if (channel ==6'b001000) nextState=ch8;
else if (channel ==6'b001001) nextState=ch9;
else if (channel ==6'b001010) nextState=ch10;
else if (channel ==6'b001011) nextState=ch11;
else if (channel ==6'b001100) nextState=ch12;
else if (channel ==6'b001101) nextState=ch13;
else if (channel ==6'b001110) nextState=ch14;
else if (channel ==6'b001111) nextState=ch15;
else if (channel ==6'b010000) nextState=ch16;
else if (channel ==6'b010001) nextState=ch17;
else if (channel ==6'b010010) nextState=ch18;
else if (channel ==6'b010011) nextState=ch19;
else if (channel ==6'b010100) nextState=ch20;
else if (channel ==6'b010101) nextState=ch21;
else if (channel ==6'b010110) nextState=ch22;
else if (channel ==6'b010111) nextState=ch23;
else if (channel ==6'b011000) nextState=ch24;
else if (channel ==6'b011001) nextState=ch25;
else if (channel ==6'b011010) nextState=ch26;
else if (channel ==6'b011011) nextState=ch27;
else if (channel ==6'b011100) nextState=ch28;
else if (channel ==6'b011101) nextState=ch29;
else if (channel ==6'b011110) nextState=ch30;
else if (channel ==6'b011111) nextState=ch31;
else if (channel ==6'b100000) nextState=ch32;
else if (channel ==6'b100001) nextState=ch33;
else if (channel ==6'b100010) nextState=ch34;
else if (channel ==6'b100011) nextState=ch35;
else if (channel ==6'b100100) nextState=ch36;
else if (channel ==6'b100101) nextState=ch37;
else if (channel ==6'b100110) nextState=ch38;
else if (channel ==6'b000000) nextState=ch0;
else if (channel ==6'b101000) nextState=ch40;
else if (channel ==6'b101001) nextState=ch41;
else if (channel ==6'b101010) nextState=ch42;
else if (channel ==6'b101011) nextState=ch43;
else if (channel ==6'b101100) nextState=ch44;
else if (channel ==6'b101101) nextState=ch45;
else if (channel ==6'b101110) nextState=ch46;
else if (channel ==6'b101111) nextState=ch47;
else if (channel ==6'b110000) nextState=ch48;
else if (channel ==6'b110001) nextState=ch49;
else if (channel ==6'b110010) nextState=ch50;
else if (channel ==6'b110011) nextState=ch51;
else if (channel ==6'b110100) nextState=ch52;
else if (channel ==6'b110101) nextState=ch53;
else if (channel ==6'b110110) nextState=ch54;
else if (channel ==6'b110111) nextState=ch55;
else if (channel ==6'b111000) nextState=ch56;
else if (channel ==6'b111001) nextState=ch57;
else if (channel ==6'b111010) nextState=ch58;
else if (channel ==6'b111011) nextState=ch59;
else if (channel ==6'b111100) nextState=ch60;
else if (channel ==6'b111101) nextState=ch61;
else if (channel ==6'b111110) nextState=ch62;
else nextState=ch63;

ch40: 
if (channel == 6'b101000) nextState=ch40;
else if (channel ==6'b000001) nextState=ch1;
else if (channel ==6'b000010) nextState=ch2;
else if (channel ==6'b000011) nextState=ch3;
else if (channel ==6'b000100) nextState=ch4;
else if (channel ==6'b000101) nextState=ch5;
else if (channel ==6'b000110) nextState=ch6;
else if (channel ==6'b000111) nextState=ch7;
else if (channel ==6'b001000) nextState=ch8;
else if (channel ==6'b001001) nextState=ch9;
else if (channel ==6'b001010) nextState=ch10;
else if (channel ==6'b001011) nextState=ch11;
else if (channel ==6'b001100) nextState=ch12;
else if (channel ==6'b001101) nextState=ch13;
else if (channel ==6'b001110) nextState=ch14;
else if (channel ==6'b001111) nextState=ch15;
else if (channel ==6'b010000) nextState=ch16;
else if (channel ==6'b010001) nextState=ch17;
else if (channel ==6'b010010) nextState=ch18;
else if (channel ==6'b010011) nextState=ch19;
else if (channel ==6'b010100) nextState=ch20;
else if (channel ==6'b010101) nextState=ch21;
else if (channel ==6'b010110) nextState=ch22;
else if (channel ==6'b010111) nextState=ch23;
else if (channel ==6'b011000) nextState=ch24;
else if (channel ==6'b011001) nextState=ch25;
else if (channel ==6'b011010) nextState=ch26;
else if (channel ==6'b011011) nextState=ch27;
else if (channel ==6'b011100) nextState=ch28;
else if (channel ==6'b011101) nextState=ch29;
else if (channel ==6'b011110) nextState=ch30;
else if (channel ==6'b011111) nextState=ch31;
else if (channel ==6'b100000) nextState=ch32;
else if (channel ==6'b100001) nextState=ch33;
else if (channel ==6'b100010) nextState=ch34;
else if (channel ==6'b100011) nextState=ch35;
else if (channel ==6'b100100) nextState=ch36;
else if (channel ==6'b100101) nextState=ch37;
else if (channel ==6'b100110) nextState=ch38;
else if (channel ==6'b100111) nextState=ch39;
else if (channel ==6'b000000) nextState=ch0;
else if (channel ==6'b101001) nextState=ch41;
else if (channel ==6'b101010) nextState=ch42;
else if (channel ==6'b101011) nextState=ch43;
else if (channel ==6'b101100) nextState=ch44;
else if (channel ==6'b101101) nextState=ch45;
else if (channel ==6'b101110) nextState=ch46;
else if (channel ==6'b101111) nextState=ch47;
else if (channel ==6'b110000) nextState=ch48;
else if (channel ==6'b110001) nextState=ch49;
else if (channel ==6'b110010) nextState=ch50;
else if (channel ==6'b110011) nextState=ch51;
else if (channel ==6'b110100) nextState=ch52;
else if (channel ==6'b110101) nextState=ch53;
else if (channel ==6'b110110) nextState=ch54;
else if (channel ==6'b110111) nextState=ch55;
else if (channel ==6'b111000) nextState=ch56;
else if (channel ==6'b111001) nextState=ch57;
else if (channel ==6'b111010) nextState=ch58;
else if (channel ==6'b111011) nextState=ch59;
else if (channel ==6'b111100) nextState=ch60;
else if (channel ==6'b111101) nextState=ch61;
else if (channel ==6'b111110) nextState=ch62;
else nextState=ch63;

ch41: 
if (channel == 6'b101001) nextState=ch41;
else if (channel ==6'b000001) nextState=ch1;
else if (channel ==6'b000010) nextState=ch2;
else if (channel ==6'b000011) nextState=ch3;
else if (channel ==6'b000100) nextState=ch4;
else if (channel ==6'b000101) nextState=ch5;
else if (channel ==6'b000110) nextState=ch6;
else if (channel ==6'b000111) nextState=ch7;
else if (channel ==6'b001000) nextState=ch8;
else if (channel ==6'b001001) nextState=ch9;
else if (channel ==6'b001010) nextState=ch10;
else if (channel ==6'b001011) nextState=ch11;
else if (channel ==6'b001100) nextState=ch12;
else if (channel ==6'b001101) nextState=ch13;
else if (channel ==6'b001110) nextState=ch14;
else if (channel ==6'b001111) nextState=ch15;
else if (channel ==6'b010000) nextState=ch16;
else if (channel ==6'b010001) nextState=ch17;
else if (channel ==6'b010010) nextState=ch18;
else if (channel ==6'b010011) nextState=ch19;
else if (channel ==6'b010100) nextState=ch20;
else if (channel ==6'b010101) nextState=ch21;
else if (channel ==6'b010110) nextState=ch22;
else if (channel ==6'b010111) nextState=ch23;
else if (channel ==6'b011000) nextState=ch24;
else if (channel ==6'b011001) nextState=ch25;
else if (channel ==6'b011010) nextState=ch26;
else if (channel ==6'b011011) nextState=ch27;
else if (channel ==6'b011100) nextState=ch28;
else if (channel ==6'b011101) nextState=ch29;
else if (channel ==6'b011110) nextState=ch30;
else if (channel ==6'b011111) nextState=ch31;
else if (channel ==6'b100000) nextState=ch32;
else if (channel ==6'b100001) nextState=ch33;
else if (channel ==6'b100010) nextState=ch34;
else if (channel ==6'b100011) nextState=ch35;
else if (channel ==6'b100100) nextState=ch36;
else if (channel ==6'b100101) nextState=ch37;
else if (channel ==6'b100110) nextState=ch38;
else if (channel ==6'b100111) nextState=ch39;
else if (channel ==6'b101000) nextState=ch40;
else if (channel ==6'b000000) nextState=ch0;
else if (channel ==6'b101010) nextState=ch42;
else if (channel ==6'b101011) nextState=ch43;
else if (channel ==6'b101100) nextState=ch44;
else if (channel ==6'b101101) nextState=ch45;
else if (channel ==6'b101110) nextState=ch46;
else if (channel ==6'b101111) nextState=ch47;
else if (channel ==6'b110000) nextState=ch48;
else if (channel ==6'b110001) nextState=ch49;
else if (channel ==6'b110010) nextState=ch50;
else if (channel ==6'b110011) nextState=ch51;
else if (channel ==6'b110100) nextState=ch52;
else if (channel ==6'b110101) nextState=ch53;
else if (channel ==6'b110110) nextState=ch54;
else if (channel ==6'b110111) nextState=ch55;
else if (channel ==6'b111000) nextState=ch56;
else if (channel ==6'b111001) nextState=ch57;
else if (channel ==6'b111010) nextState=ch58;
else if (channel ==6'b111011) nextState=ch59;
else if (channel ==6'b111100) nextState=ch60;
else if (channel ==6'b111101) nextState=ch61;
else if (channel ==6'b111110) nextState=ch62;
else nextState=ch63;

ch42: 
if (channel == 6'b101010) nextState=ch42;
else if (channel ==6'b000001) nextState=ch1;
else if (channel ==6'b000010) nextState=ch2;
else if (channel ==6'b000011) nextState=ch3;
else if (channel ==6'b000100) nextState=ch4;
else if (channel ==6'b000101) nextState=ch5;
else if (channel ==6'b000110) nextState=ch6;
else if (channel ==6'b000111) nextState=ch7;
else if (channel ==6'b001000) nextState=ch8;
else if (channel ==6'b001001) nextState=ch9;
else if (channel ==6'b001010) nextState=ch10;
else if (channel ==6'b001011) nextState=ch11;
else if (channel ==6'b001100) nextState=ch12;
else if (channel ==6'b001101) nextState=ch13;
else if (channel ==6'b001110) nextState=ch14;
else if (channel ==6'b001111) nextState=ch15;
else if (channel ==6'b010000) nextState=ch16;
else if (channel ==6'b010001) nextState=ch17;
else if (channel ==6'b010010) nextState=ch18;
else if (channel ==6'b010011) nextState=ch19;
else if (channel ==6'b010100) nextState=ch20;
else if (channel ==6'b010101) nextState=ch21;
else if (channel ==6'b010110) nextState=ch22;
else if (channel ==6'b010111) nextState=ch23;
else if (channel ==6'b011000) nextState=ch24;
else if (channel ==6'b011001) nextState=ch25;
else if (channel ==6'b011010) nextState=ch26;
else if (channel ==6'b011011) nextState=ch27;
else if (channel ==6'b011100) nextState=ch28;
else if (channel ==6'b011101) nextState=ch29;
else if (channel ==6'b011110) nextState=ch30;
else if (channel ==6'b011111) nextState=ch31;
else if (channel ==6'b100000) nextState=ch32;
else if (channel ==6'b100001) nextState=ch33;
else if (channel ==6'b100010) nextState=ch34;
else if (channel ==6'b100011) nextState=ch35;
else if (channel ==6'b100100) nextState=ch36;
else if (channel ==6'b100101) nextState=ch37;
else if (channel ==6'b100110) nextState=ch38;
else if (channel ==6'b100111) nextState=ch39;
else if (channel ==6'b101000) nextState=ch40;
else if (channel ==6'b101001) nextState=ch41;
else if (channel ==6'b000000) nextState=ch0;
else if (channel ==6'b101011) nextState=ch43;
else if (channel ==6'b101100) nextState=ch44;
else if (channel ==6'b101101) nextState=ch45;
else if (channel ==6'b101110) nextState=ch46;
else if (channel ==6'b101111) nextState=ch47;
else if (channel ==6'b110000) nextState=ch48;
else if (channel ==6'b110001) nextState=ch49;
else if (channel ==6'b110010) nextState=ch50;
else if (channel ==6'b110011) nextState=ch51;
else if (channel ==6'b110100) nextState=ch52;
else if (channel ==6'b110101) nextState=ch53;
else if (channel ==6'b110110) nextState=ch54;
else if (channel ==6'b110111) nextState=ch55;
else if (channel ==6'b111000) nextState=ch56;
else if (channel ==6'b111001) nextState=ch57;
else if (channel ==6'b111010) nextState=ch58;
else if (channel ==6'b111011) nextState=ch59;
else if (channel ==6'b111100) nextState=ch60;
else if (channel ==6'b111101) nextState=ch61;
else if (channel ==6'b111110) nextState=ch62;
else nextState=ch63;

ch43: 
if (channel == 6'b101011) nextState=ch43;
else if (channel ==6'b000001) nextState=ch1;
else if (channel ==6'b000010) nextState=ch2;
else if (channel ==6'b000011) nextState=ch3;
else if (channel ==6'b000100) nextState=ch4;
else if (channel ==6'b000101) nextState=ch5;
else if (channel ==6'b000110) nextState=ch6;
else if (channel ==6'b000111) nextState=ch7;
else if (channel ==6'b001000) nextState=ch8;
else if (channel ==6'b001001) nextState=ch9;
else if (channel ==6'b001010) nextState=ch10;
else if (channel ==6'b001011) nextState=ch11;
else if (channel ==6'b001100) nextState=ch12;
else if (channel ==6'b001101) nextState=ch13;
else if (channel ==6'b001110) nextState=ch14;
else if (channel ==6'b001111) nextState=ch15;
else if (channel ==6'b010000) nextState=ch16;
else if (channel ==6'b010001) nextState=ch17;
else if (channel ==6'b010010) nextState=ch18;
else if (channel ==6'b010011) nextState=ch19;
else if (channel ==6'b010100) nextState=ch20;
else if (channel ==6'b010101) nextState=ch21;
else if (channel ==6'b010110) nextState=ch22;
else if (channel ==6'b010111) nextState=ch23;
else if (channel ==6'b011000) nextState=ch24;
else if (channel ==6'b011001) nextState=ch25;
else if (channel ==6'b011010) nextState=ch26;
else if (channel ==6'b011011) nextState=ch27;
else if (channel ==6'b011100) nextState=ch28;
else if (channel ==6'b011101) nextState=ch29;
else if (channel ==6'b011110) nextState=ch30;
else if (channel ==6'b011111) nextState=ch31;
else if (channel ==6'b100000) nextState=ch32;
else if (channel ==6'b100001) nextState=ch33;
else if (channel ==6'b100010) nextState=ch34;
else if (channel ==6'b100011) nextState=ch35;
else if (channel ==6'b100100) nextState=ch36;
else if (channel ==6'b100101) nextState=ch37;
else if (channel ==6'b100110) nextState=ch38;
else if (channel ==6'b100111) nextState=ch39;
else if (channel ==6'b101000) nextState=ch40;
else if (channel ==6'b101001) nextState=ch41;
else if (channel ==6'b101010) nextState=ch42;
else if (channel ==6'b000000) nextState=ch0;
else if (channel ==6'b101100) nextState=ch44;
else if (channel ==6'b101101) nextState=ch45;
else if (channel ==6'b101110) nextState=ch46;
else if (channel ==6'b101111) nextState=ch47;
else if (channel ==6'b110000) nextState=ch48;
else if (channel ==6'b110001) nextState=ch49;
else if (channel ==6'b110010) nextState=ch50;
else if (channel ==6'b110011) nextState=ch51;
else if (channel ==6'b110100) nextState=ch52;
else if (channel ==6'b110101) nextState=ch53;
else if (channel ==6'b110110) nextState=ch54;
else if (channel ==6'b110111) nextState=ch55;
else if (channel ==6'b111000) nextState=ch56;
else if (channel ==6'b111001) nextState=ch57;
else if (channel ==6'b111010) nextState=ch58;
else if (channel ==6'b111011) nextState=ch59;
else if (channel ==6'b111100) nextState=ch60;
else if (channel ==6'b111101) nextState=ch61;
else if (channel ==6'b111110) nextState=ch62;
else nextState=ch63;

ch44: 
if (channel == 6'b101100) nextState=ch44;
else if (channel ==6'b000001) nextState=ch1;
else if (channel ==6'b000010) nextState=ch2;
else if (channel ==6'b000011) nextState=ch3;
else if (channel ==6'b000100) nextState=ch4;
else if (channel ==6'b000101) nextState=ch5;
else if (channel ==6'b000110) nextState=ch6;
else if (channel ==6'b000111) nextState=ch7;
else if (channel ==6'b001000) nextState=ch8;
else if (channel ==6'b001001) nextState=ch9;
else if (channel ==6'b001010) nextState=ch10;
else if (channel ==6'b001011) nextState=ch11;
else if (channel ==6'b001100) nextState=ch12;
else if (channel ==6'b001101) nextState=ch13;
else if (channel ==6'b001110) nextState=ch14;
else if (channel ==6'b001111) nextState=ch15;
else if (channel ==6'b010000) nextState=ch16;
else if (channel ==6'b010001) nextState=ch17;
else if (channel ==6'b010010) nextState=ch18;
else if (channel ==6'b010011) nextState=ch19;
else if (channel ==6'b010100) nextState=ch20;
else if (channel ==6'b010101) nextState=ch21;
else if (channel ==6'b010110) nextState=ch22;
else if (channel ==6'b010111) nextState=ch23;
else if (channel ==6'b011000) nextState=ch24;
else if (channel ==6'b011001) nextState=ch25;
else if (channel ==6'b011010) nextState=ch26;
else if (channel ==6'b011011) nextState=ch27;
else if (channel ==6'b011100) nextState=ch28;
else if (channel ==6'b011101) nextState=ch29;
else if (channel ==6'b011110) nextState=ch30;
else if (channel ==6'b011111) nextState=ch31;
else if (channel ==6'b100000) nextState=ch32;
else if (channel ==6'b100001) nextState=ch33;
else if (channel ==6'b100010) nextState=ch34;
else if (channel ==6'b100011) nextState=ch35;
else if (channel ==6'b100100) nextState=ch36;
else if (channel ==6'b100101) nextState=ch37;
else if (channel ==6'b100110) nextState=ch38;
else if (channel ==6'b100111) nextState=ch39;
else if (channel ==6'b101000) nextState=ch40;
else if (channel ==6'b101001) nextState=ch41;
else if (channel ==6'b101010) nextState=ch42;
else if (channel ==6'b101011) nextState=ch43;
else if (channel ==6'b000000) nextState=ch0;
else if (channel ==6'b101101) nextState=ch45;
else if (channel ==6'b101110) nextState=ch46;
else if (channel ==6'b101111) nextState=ch47;
else if (channel ==6'b110000) nextState=ch48;
else if (channel ==6'b110001) nextState=ch49;
else if (channel ==6'b110010) nextState=ch50;
else if (channel ==6'b110011) nextState=ch51;
else if (channel ==6'b110100) nextState=ch52;
else if (channel ==6'b110101) nextState=ch53;
else if (channel ==6'b110110) nextState=ch54;
else if (channel ==6'b110111) nextState=ch55;
else if (channel ==6'b111000) nextState=ch56;
else if (channel ==6'b111001) nextState=ch57;
else if (channel ==6'b111010) nextState=ch58;
else if (channel ==6'b111011) nextState=ch59;
else if (channel ==6'b111100) nextState=ch60;
else if (channel ==6'b111101) nextState=ch61;
else if (channel ==6'b111110) nextState=ch62;
else nextState=ch63;

ch45: 
if (channel == 6'b101101) nextState=ch45;
else if (channel ==6'b000001) nextState=ch1;
else if (channel ==6'b000010) nextState=ch2;
else if (channel ==6'b000011) nextState=ch3;
else if (channel ==6'b000100) nextState=ch4;
else if (channel ==6'b000101) nextState=ch5;
else if (channel ==6'b000110) nextState=ch6;
else if (channel ==6'b000111) nextState=ch7;
else if (channel ==6'b001000) nextState=ch8;
else if (channel ==6'b001001) nextState=ch9;
else if (channel ==6'b001010) nextState=ch10;
else if (channel ==6'b001011) nextState=ch11;
else if (channel ==6'b001100) nextState=ch12;
else if (channel ==6'b001101) nextState=ch13;
else if (channel ==6'b001110) nextState=ch14;
else if (channel ==6'b001111) nextState=ch15;
else if (channel ==6'b010000) nextState=ch16;
else if (channel ==6'b010001) nextState=ch17;
else if (channel ==6'b010010) nextState=ch18;
else if (channel ==6'b010011) nextState=ch19;
else if (channel ==6'b010100) nextState=ch20;
else if (channel ==6'b010101) nextState=ch21;
else if (channel ==6'b010110) nextState=ch22;
else if (channel ==6'b010111) nextState=ch23;
else if (channel ==6'b011000) nextState=ch24;
else if (channel ==6'b011001) nextState=ch25;
else if (channel ==6'b011010) nextState=ch26;
else if (channel ==6'b011011) nextState=ch27;
else if (channel ==6'b011100) nextState=ch28;
else if (channel ==6'b011101) nextState=ch29;
else if (channel ==6'b011110) nextState=ch30;
else if (channel ==6'b011111) nextState=ch31;
else if (channel ==6'b100000) nextState=ch32;
else if (channel ==6'b100001) nextState=ch33;
else if (channel ==6'b100010) nextState=ch34;
else if (channel ==6'b100011) nextState=ch35;
else if (channel ==6'b100100) nextState=ch36;
else if (channel ==6'b100101) nextState=ch37;
else if (channel ==6'b100110) nextState=ch38;
else if (channel ==6'b100111) nextState=ch39;
else if (channel ==6'b101000) nextState=ch40;
else if (channel ==6'b101001) nextState=ch41;
else if (channel ==6'b101010) nextState=ch42;
else if (channel ==6'b101011) nextState=ch43;
else if (channel ==6'b101100) nextState=ch44;
else if (channel ==6'b000000) nextState=ch45;
else if (channel ==6'b101110) nextState=ch46;
else if (channel ==6'b101111) nextState=ch47;
else if (channel ==6'b110000) nextState=ch48;
else if (channel ==6'b110001) nextState=ch49;
else if (channel ==6'b110010) nextState=ch50;
else if (channel ==6'b110011) nextState=ch51;
else if (channel ==6'b110100) nextState=ch52;
else if (channel ==6'b110101) nextState=ch53;
else if (channel ==6'b110110) nextState=ch54;
else if (channel ==6'b110111) nextState=ch55;
else if (channel ==6'b111000) nextState=ch56;
else if (channel ==6'b111001) nextState=ch57;
else if (channel ==6'b111010) nextState=ch58;
else if (channel ==6'b111011) nextState=ch59;
else if (channel ==6'b111100) nextState=ch60;
else if (channel ==6'b111101) nextState=ch61;
else if (channel ==6'b111110) nextState=ch62;
else nextState=ch63;

ch46: 
if (channel == 6'b101110) nextState=ch46;
else if (channel ==6'b000001) nextState=ch1;
else if (channel ==6'b000010) nextState=ch2;
else if (channel ==6'b000011) nextState=ch3;
else if (channel ==6'b000100) nextState=ch4;
else if (channel ==6'b000101) nextState=ch5;
else if (channel ==6'b000110) nextState=ch6;
else if (channel ==6'b000111) nextState=ch7;
else if (channel ==6'b001000) nextState=ch8;
else if (channel ==6'b001001) nextState=ch9;
else if (channel ==6'b001010) nextState=ch10;
else if (channel ==6'b001011) nextState=ch11;
else if (channel ==6'b001100) nextState=ch12;
else if (channel ==6'b001101) nextState=ch13;
else if (channel ==6'b001110) nextState=ch14;
else if (channel ==6'b001111) nextState=ch15;
else if (channel ==6'b010000) nextState=ch16;
else if (channel ==6'b010001) nextState=ch17;
else if (channel ==6'b010010) nextState=ch18;
else if (channel ==6'b010011) nextState=ch19;
else if (channel ==6'b010100) nextState=ch20;
else if (channel ==6'b010101) nextState=ch21;
else if (channel ==6'b010110) nextState=ch22;
else if (channel ==6'b010111) nextState=ch23;
else if (channel ==6'b011000) nextState=ch24;
else if (channel ==6'b011001) nextState=ch25;
else if (channel ==6'b011010) nextState=ch26;
else if (channel ==6'b011011) nextState=ch27;
else if (channel ==6'b011100) nextState=ch28;
else if (channel ==6'b011101) nextState=ch29;
else if (channel ==6'b011110) nextState=ch30;
else if (channel ==6'b011111) nextState=ch31;
else if (channel ==6'b100000) nextState=ch32;
else if (channel ==6'b100001) nextState=ch33;
else if (channel ==6'b100010) nextState=ch34;
else if (channel ==6'b100011) nextState=ch35;
else if (channel ==6'b100100) nextState=ch36;
else if (channel ==6'b100101) nextState=ch37;
else if (channel ==6'b100110) nextState=ch38;
else if (channel ==6'b100111) nextState=ch39;
else if (channel ==6'b101000) nextState=ch40;
else if (channel ==6'b101001) nextState=ch41;
else if (channel ==6'b101010) nextState=ch42;
else if (channel ==6'b101011) nextState=ch43;
else if (channel ==6'b101100) nextState=ch44;
else if (channel ==6'b101101) nextState=ch45;
else if (channel ==6'b000000) nextState=ch0;
else if (channel ==6'b101111) nextState=ch47;
else if (channel ==6'b110000) nextState=ch48;
else if (channel ==6'b110001) nextState=ch49;
else if (channel ==6'b110010) nextState=ch50;
else if (channel ==6'b110011) nextState=ch51;
else if (channel ==6'b110100) nextState=ch52;
else if (channel ==6'b110101) nextState=ch53;
else if (channel ==6'b110110) nextState=ch54;
else if (channel ==6'b110111) nextState=ch55;
else if (channel ==6'b111000) nextState=ch56;
else if (channel ==6'b111001) nextState=ch57;
else if (channel ==6'b111010) nextState=ch58;
else if (channel ==6'b111011) nextState=ch59;
else if (channel ==6'b111100) nextState=ch60;
else if (channel ==6'b111101) nextState=ch61;
else if (channel ==6'b111110) nextState=ch62;
else nextState=ch63;

ch47: 
if (channel == 6'b101111) nextState=ch47;
else if (channel ==6'b000001) nextState=ch1;
else if (channel ==6'b000010) nextState=ch2;
else if (channel ==6'b000011) nextState=ch3;
else if (channel ==6'b000100) nextState=ch4;
else if (channel ==6'b000101) nextState=ch5;
else if (channel ==6'b000110) nextState=ch6;
else if (channel ==6'b000111) nextState=ch7;
else if (channel ==6'b001000) nextState=ch8;
else if (channel ==6'b001001) nextState=ch9;
else if (channel ==6'b001010) nextState=ch10;
else if (channel ==6'b001011) nextState=ch11;
else if (channel ==6'b001100) nextState=ch12;
else if (channel ==6'b001101) nextState=ch13;
else if (channel ==6'b001110) nextState=ch14;
else if (channel ==6'b001111) nextState=ch15;
else if (channel ==6'b010000) nextState=ch16;
else if (channel ==6'b010001) nextState=ch17;
else if (channel ==6'b010010) nextState=ch18;
else if (channel ==6'b010011) nextState=ch19;
else if (channel ==6'b010100) nextState=ch20;
else if (channel ==6'b010101) nextState=ch21;
else if (channel ==6'b010110) nextState=ch22;
else if (channel ==6'b010111) nextState=ch23;
else if (channel ==6'b011000) nextState=ch24;
else if (channel ==6'b011001) nextState=ch25;
else if (channel ==6'b011010) nextState=ch26;
else if (channel ==6'b011011) nextState=ch27;
else if (channel ==6'b011100) nextState=ch28;
else if (channel ==6'b011101) nextState=ch29;
else if (channel ==6'b011110) nextState=ch30;
else if (channel ==6'b011111) nextState=ch31;
else if (channel ==6'b100000) nextState=ch32;
else if (channel ==6'b100001) nextState=ch33;
else if (channel ==6'b100010) nextState=ch34;
else if (channel ==6'b100011) nextState=ch35;
else if (channel ==6'b100100) nextState=ch36;
else if (channel ==6'b100101) nextState=ch37;
else if (channel ==6'b100110) nextState=ch38;
else if (channel ==6'b100111) nextState=ch39;
else if (channel ==6'b101000) nextState=ch40;
else if (channel ==6'b101001) nextState=ch41;
else if (channel ==6'b101010) nextState=ch42;
else if (channel ==6'b101011) nextState=ch43;
else if (channel ==6'b101100) nextState=ch44;
else if (channel ==6'b101101) nextState=ch45;
else if (channel ==6'b101110) nextState=ch46;
else if (channel ==6'b000000) nextState=ch0;
else if (channel ==6'b110000) nextState=ch48;
else if (channel ==6'b110001) nextState=ch49;
else if (channel ==6'b110010) nextState=ch50;
else if (channel ==6'b110011) nextState=ch51;
else if (channel ==6'b110100) nextState=ch52;
else if (channel ==6'b110101) nextState=ch53;
else if (channel ==6'b110110) nextState=ch54;
else if (channel ==6'b110111) nextState=ch55;
else if (channel ==6'b111000) nextState=ch56;
else if (channel ==6'b111001) nextState=ch57;
else if (channel ==6'b111010) nextState=ch58;
else if (channel ==6'b111011) nextState=ch59;
else if (channel ==6'b111100) nextState=ch60;
else if (channel ==6'b111101) nextState=ch61;
else if (channel ==6'b111110) nextState=ch62;
else nextState=ch63;

ch48: 
if (channel == 6'b110000) nextState=ch48;
else if (channel ==6'b000001) nextState=ch1;
else if (channel ==6'b000010) nextState=ch2;
else if (channel ==6'b000011) nextState=ch3;
else if (channel ==6'b000100) nextState=ch4;
else if (channel ==6'b000101) nextState=ch5;
else if (channel ==6'b000110) nextState=ch6;
else if (channel ==6'b000111) nextState=ch7;
else if (channel ==6'b001000) nextState=ch8;
else if (channel ==6'b001001) nextState=ch9;
else if (channel ==6'b001010) nextState=ch10;
else if (channel ==6'b001011) nextState=ch11;
else if (channel ==6'b001100) nextState=ch12;
else if (channel ==6'b001101) nextState=ch13;
else if (channel ==6'b001110) nextState=ch14;
else if (channel ==6'b001111) nextState=ch15;
else if (channel ==6'b010000) nextState=ch16;
else if (channel ==6'b010001) nextState=ch17;
else if (channel ==6'b010010) nextState=ch18;
else if (channel ==6'b010011) nextState=ch19;
else if (channel ==6'b010100) nextState=ch20;
else if (channel ==6'b010101) nextState=ch21;
else if (channel ==6'b010110) nextState=ch22;
else if (channel ==6'b010111) nextState=ch23;
else if (channel ==6'b011000) nextState=ch24;
else if (channel ==6'b011001) nextState=ch25;
else if (channel ==6'b011010) nextState=ch26;
else if (channel ==6'b011011) nextState=ch27;
else if (channel ==6'b011100) nextState=ch28;
else if (channel ==6'b011101) nextState=ch29;
else if (channel ==6'b011110) nextState=ch30;
else if (channel ==6'b011111) nextState=ch31;
else if (channel ==6'b100000) nextState=ch32;
else if (channel ==6'b100001) nextState=ch33;
else if (channel ==6'b100010) nextState=ch34;
else if (channel ==6'b100011) nextState=ch35;
else if (channel ==6'b100100) nextState=ch36;
else if (channel ==6'b100101) nextState=ch37;
else if (channel ==6'b100110) nextState=ch38;
else if (channel ==6'b100111) nextState=ch39;
else if (channel ==6'b101000) nextState=ch40;
else if (channel ==6'b101001) nextState=ch41;
else if (channel ==6'b101010) nextState=ch42;
else if (channel ==6'b101011) nextState=ch43;
else if (channel ==6'b101100) nextState=ch44;
else if (channel ==6'b101101) nextState=ch45;
else if (channel ==6'b101110) nextState=ch46;
else if (channel ==6'b101111) nextState=ch47;
else if (channel ==6'b000000) nextState=ch0;
else if (channel ==6'b110001) nextState=ch49;
else if (channel ==6'b110010) nextState=ch50;
else if (channel ==6'b110011) nextState=ch51;
else if (channel ==6'b110100) nextState=ch52;
else if (channel ==6'b110101) nextState=ch53;
else if (channel ==6'b110110) nextState=ch54;
else if (channel ==6'b110111) nextState=ch55;
else if (channel ==6'b111000) nextState=ch56;
else if (channel ==6'b111001) nextState=ch57;
else if (channel ==6'b111010) nextState=ch58;
else if (channel ==6'b111011) nextState=ch59;
else if (channel ==6'b111100) nextState=ch60;
else if (channel ==6'b111101) nextState=ch61;
else if (channel ==6'b111110) nextState=ch62;
else nextState=ch63;

ch49: 
if (channel == 6'b110001) nextState=ch49;
else if (channel ==6'b000001) nextState=ch1;
else if (channel ==6'b000010) nextState=ch2;
else if (channel ==6'b000011) nextState=ch3;
else if (channel ==6'b000100) nextState=ch4;
else if (channel ==6'b000101) nextState=ch5;
else if (channel ==6'b000110) nextState=ch6;
else if (channel ==6'b000111) nextState=ch7;
else if (channel ==6'b001000) nextState=ch8;
else if (channel ==6'b001001) nextState=ch9;
else if (channel ==6'b001010) nextState=ch10;
else if (channel ==6'b001011) nextState=ch11;
else if (channel ==6'b001100) nextState=ch12;
else if (channel ==6'b001101) nextState=ch13;
else if (channel ==6'b001110) nextState=ch14;
else if (channel ==6'b001111) nextState=ch15;
else if (channel ==6'b010000) nextState=ch16;
else if (channel ==6'b010001) nextState=ch17;
else if (channel ==6'b010010) nextState=ch18;
else if (channel ==6'b010011) nextState=ch19;
else if (channel ==6'b010100) nextState=ch20;
else if (channel ==6'b010101) nextState=ch21;
else if (channel ==6'b010110) nextState=ch22;
else if (channel ==6'b010111) nextState=ch23;
else if (channel ==6'b011000) nextState=ch24;
else if (channel ==6'b011001) nextState=ch25;
else if (channel ==6'b011010) nextState=ch26;
else if (channel ==6'b011011) nextState=ch27;
else if (channel ==6'b011100) nextState=ch28;
else if (channel ==6'b011101) nextState=ch29;
else if (channel ==6'b011110) nextState=ch30;
else if (channel ==6'b011111) nextState=ch31;
else if (channel ==6'b100000) nextState=ch32;
else if (channel ==6'b100001) nextState=ch33;
else if (channel ==6'b100010) nextState=ch34;
else if (channel ==6'b100011) nextState=ch35;
else if (channel ==6'b100100) nextState=ch36;
else if (channel ==6'b100101) nextState=ch37;
else if (channel ==6'b100110) nextState=ch38;
else if (channel ==6'b100111) nextState=ch39;
else if (channel ==6'b101000) nextState=ch40;
else if (channel ==6'b101001) nextState=ch41;
else if (channel ==6'b101010) nextState=ch42;
else if (channel ==6'b101011) nextState=ch43;
else if (channel ==6'b101100) nextState=ch44;
else if (channel ==6'b101101) nextState=ch45;
else if (channel ==6'b101110) nextState=ch46;
else if (channel ==6'b101111) nextState=ch47;
else if (channel ==6'b110000) nextState=ch48;
else if (channel ==6'b000000) nextState=ch0;
else if (channel ==6'b110010) nextState=ch50;
else if (channel ==6'b110011) nextState=ch51;
else if (channel ==6'b110100) nextState=ch52;
else if (channel ==6'b110101) nextState=ch53;
else if (channel ==6'b110110) nextState=ch54;
else if (channel ==6'b110111) nextState=ch55;
else if (channel ==6'b111000) nextState=ch56;
else if (channel ==6'b111001) nextState=ch57;
else if (channel ==6'b111010) nextState=ch58;
else if (channel ==6'b111011) nextState=ch59;
else if (channel ==6'b111100) nextState=ch60;
else if (channel ==6'b111101) nextState=ch61;
else if (channel ==6'b111110) nextState=ch62;
else nextState=ch63;

ch50: 
if (channel == 6'b110010) nextState=ch50;
else if (channel ==6'b000001) nextState=ch1;
else if (channel ==6'b000010) nextState=ch2;
else if (channel ==6'b000011) nextState=ch3;
else if (channel ==6'b000100) nextState=ch4;
else if (channel ==6'b000101) nextState=ch5;
else if (channel ==6'b000110) nextState=ch6;
else if (channel ==6'b000111) nextState=ch7;
else if (channel ==6'b001000) nextState=ch8;
else if (channel ==6'b001001) nextState=ch9;
else if (channel ==6'b001010) nextState=ch10;
else if (channel ==6'b001011) nextState=ch11;
else if (channel ==6'b001100) nextState=ch12;
else if (channel ==6'b001101) nextState=ch13;
else if (channel ==6'b001110) nextState=ch14;
else if (channel ==6'b001111) nextState=ch15;
else if (channel ==6'b010000) nextState=ch16;
else if (channel ==6'b010001) nextState=ch17;
else if (channel ==6'b010010) nextState=ch18;
else if (channel ==6'b010011) nextState=ch19;
else if (channel ==6'b010100) nextState=ch20;
else if (channel ==6'b010101) nextState=ch21;
else if (channel ==6'b010110) nextState=ch22;
else if (channel ==6'b010111) nextState=ch23;
else if (channel ==6'b011000) nextState=ch24;
else if (channel ==6'b011001) nextState=ch25;
else if (channel ==6'b011010) nextState=ch26;
else if (channel ==6'b011011) nextState=ch27;
else if (channel ==6'b011100) nextState=ch28;
else if (channel ==6'b011101) nextState=ch29;
else if (channel ==6'b011110) nextState=ch30;
else if (channel ==6'b011111) nextState=ch31;
else if (channel ==6'b100000) nextState=ch32;
else if (channel ==6'b100001) nextState=ch33;
else if (channel ==6'b100010) nextState=ch34;
else if (channel ==6'b100011) nextState=ch35;
else if (channel ==6'b100100) nextState=ch36;
else if (channel ==6'b100101) nextState=ch37;
else if (channel ==6'b100110) nextState=ch38;
else if (channel ==6'b100111) nextState=ch39;
else if (channel ==6'b101000) nextState=ch40;
else if (channel ==6'b101001) nextState=ch41;
else if (channel ==6'b101010) nextState=ch42;
else if (channel ==6'b101011) nextState=ch43;
else if (channel ==6'b101100) nextState=ch44;
else if (channel ==6'b101101) nextState=ch45;
else if (channel ==6'b101110) nextState=ch46;
else if (channel ==6'b101111) nextState=ch47;
else if (channel ==6'b110000) nextState=ch48;
else if (channel ==6'b110001) nextState=ch49;
else if (channel ==6'b000000) nextState=ch0;
else if (channel ==6'b110011) nextState=ch51;
else if (channel ==6'b110100) nextState=ch52;
else if (channel ==6'b110101) nextState=ch53;
else if (channel ==6'b110110) nextState=ch54;
else if (channel ==6'b110111) nextState=ch55;
else if (channel ==6'b111000) nextState=ch56;
else if (channel ==6'b111001) nextState=ch57;
else if (channel ==6'b111010) nextState=ch58;
else if (channel ==6'b111011) nextState=ch59;
else if (channel ==6'b111100) nextState=ch60;
else if (channel ==6'b111101) nextState=ch61;
else if (channel ==6'b111110) nextState=ch62;
else nextState=ch63;

ch51: 
if (channel == 6'b110011) nextState=ch51;
else if (channel ==6'b000001) nextState=ch1;
else if (channel ==6'b000010) nextState=ch2;
else if (channel ==6'b000011) nextState=ch3;
else if (channel ==6'b000100) nextState=ch4;
else if (channel ==6'b000101) nextState=ch5;
else if (channel ==6'b000110) nextState=ch6;
else if (channel ==6'b000111) nextState=ch7;
else if (channel ==6'b001000) nextState=ch8;
else if (channel ==6'b001001) nextState=ch9;
else if (channel ==6'b001010) nextState=ch10;
else if (channel ==6'b001011) nextState=ch11;
else if (channel ==6'b001100) nextState=ch12;
else if (channel ==6'b001101) nextState=ch13;
else if (channel ==6'b001110) nextState=ch14;
else if (channel ==6'b001111) nextState=ch15;
else if (channel ==6'b010000) nextState=ch16;
else if (channel ==6'b010001) nextState=ch17;
else if (channel ==6'b010010) nextState=ch18;
else if (channel ==6'b010011) nextState=ch19;
else if (channel ==6'b010100) nextState=ch20;
else if (channel ==6'b010101) nextState=ch21;
else if (channel ==6'b010110) nextState=ch22;
else if (channel ==6'b010111) nextState=ch23;
else if (channel ==6'b011000) nextState=ch24;
else if (channel ==6'b011001) nextState=ch25;
else if (channel ==6'b011010) nextState=ch26;
else if (channel ==6'b011011) nextState=ch27;
else if (channel ==6'b011100) nextState=ch28;
else if (channel ==6'b011101) nextState=ch29;
else if (channel ==6'b011110) nextState=ch30;
else if (channel ==6'b011111) nextState=ch31;
else if (channel ==6'b100000) nextState=ch32;
else if (channel ==6'b100001) nextState=ch33;
else if (channel ==6'b100010) nextState=ch34;
else if (channel ==6'b100011) nextState=ch35;
else if (channel ==6'b100100) nextState=ch36;
else if (channel ==6'b100101) nextState=ch37;
else if (channel ==6'b100110) nextState=ch38;
else if (channel ==6'b100111) nextState=ch39;
else if (channel ==6'b101000) nextState=ch40;
else if (channel ==6'b101001) nextState=ch41;
else if (channel ==6'b101010) nextState=ch42;
else if (channel ==6'b101011) nextState=ch43;
else if (channel ==6'b101100) nextState=ch44;
else if (channel ==6'b101101) nextState=ch45;
else if (channel ==6'b101110) nextState=ch46;
else if (channel ==6'b101111) nextState=ch47;
else if (channel ==6'b110000) nextState=ch48;
else if (channel ==6'b110001) nextState=ch49;
else if (channel ==6'b110010) nextState=ch50;
else if (channel ==6'b000000) nextState=ch0;
else if (channel ==6'b110100) nextState=ch52;
else if (channel ==6'b110101) nextState=ch53;
else if (channel ==6'b110110) nextState=ch54;
else if (channel ==6'b110111) nextState=ch55;
else if (channel ==6'b111000) nextState=ch56;
else if (channel ==6'b111001) nextState=ch57;
else if (channel ==6'b111010) nextState=ch58;
else if (channel ==6'b111011) nextState=ch59;
else if (channel ==6'b111100) nextState=ch60;
else if (channel ==6'b111101) nextState=ch61;
else if (channel ==6'b111110) nextState=ch62;
else nextState=ch63;

ch52: 
if (channel == 6'b110100) nextState=ch52;
else if (channel ==6'b000001) nextState=ch1;
else if (channel ==6'b000010) nextState=ch2;
else if (channel ==6'b000011) nextState=ch3;
else if (channel ==6'b000100) nextState=ch4;
else if (channel ==6'b000101) nextState=ch5;
else if (channel ==6'b000110) nextState=ch6;
else if (channel ==6'b000111) nextState=ch7;
else if (channel ==6'b001000) nextState=ch8;
else if (channel ==6'b001001) nextState=ch9;
else if (channel ==6'b001010) nextState=ch10;
else if (channel ==6'b001011) nextState=ch11;
else if (channel ==6'b001100) nextState=ch12;
else if (channel ==6'b001101) nextState=ch13;
else if (channel ==6'b001110) nextState=ch14;
else if (channel ==6'b001111) nextState=ch15;
else if (channel ==6'b010000) nextState=ch16;
else if (channel ==6'b010001) nextState=ch17;
else if (channel ==6'b010010) nextState=ch18;
else if (channel ==6'b010011) nextState=ch19;
else if (channel ==6'b010100) nextState=ch20;
else if (channel ==6'b010101) nextState=ch21;
else if (channel ==6'b010110) nextState=ch22;
else if (channel ==6'b010111) nextState=ch23;
else if (channel ==6'b011000) nextState=ch24;
else if (channel ==6'b011001) nextState=ch25;
else if (channel ==6'b011010) nextState=ch26;
else if (channel ==6'b011011) nextState=ch27;
else if (channel ==6'b011100) nextState=ch28;
else if (channel ==6'b011101) nextState=ch29;
else if (channel ==6'b011110) nextState=ch30;
else if (channel ==6'b011111) nextState=ch31;
else if (channel ==6'b100000) nextState=ch32;
else if (channel ==6'b100001) nextState=ch33;
else if (channel ==6'b100010) nextState=ch34;
else if (channel ==6'b100011) nextState=ch35;
else if (channel ==6'b100100) nextState=ch36;
else if (channel ==6'b100101) nextState=ch37;
else if (channel ==6'b100110) nextState=ch38;
else if (channel ==6'b100111) nextState=ch39;
else if (channel ==6'b101000) nextState=ch40;
else if (channel ==6'b101001) nextState=ch41;
else if (channel ==6'b101010) nextState=ch42;
else if (channel ==6'b101011) nextState=ch43;
else if (channel ==6'b101100) nextState=ch44;
else if (channel ==6'b101101) nextState=ch45;
else if (channel ==6'b101110) nextState=ch46;
else if (channel ==6'b101111) nextState=ch47;
else if (channel ==6'b110000) nextState=ch48;
else if (channel ==6'b110001) nextState=ch49;
else if (channel ==6'b110010) nextState=ch50;
else if (channel ==6'b110011) nextState=ch51;
else if (channel ==6'b000000) nextState=ch0;
else if (channel ==6'b110101) nextState=ch53;
else if (channel ==6'b110110) nextState=ch54;
else if (channel ==6'b110111) nextState=ch55;
else if (channel ==6'b111000) nextState=ch56;
else if (channel ==6'b111001) nextState=ch57;
else if (channel ==6'b111010) nextState=ch58;
else if (channel ==6'b111011) nextState=ch59;
else if (channel ==6'b111100) nextState=ch60;
else if (channel ==6'b111101) nextState=ch61;
else if (channel ==6'b111110) nextState=ch62;
else nextState=ch63;

ch53: 
if (channel == 6'b110101) nextState=ch53;
else if (channel ==6'b000001) nextState=ch1;
else if (channel ==6'b000010) nextState=ch2;
else if (channel ==6'b000011) nextState=ch3;
else if (channel ==6'b000100) nextState=ch4;
else if (channel ==6'b000101) nextState=ch5;
else if (channel ==6'b000110) nextState=ch6;
else if (channel ==6'b000111) nextState=ch7;
else if (channel ==6'b001000) nextState=ch8;
else if (channel ==6'b001001) nextState=ch9;
else if (channel ==6'b001010) nextState=ch10;
else if (channel ==6'b001011) nextState=ch11;
else if (channel ==6'b001100) nextState=ch12;
else if (channel ==6'b001101) nextState=ch13;
else if (channel ==6'b001110) nextState=ch14;
else if (channel ==6'b001111) nextState=ch15;
else if (channel ==6'b010000) nextState=ch16;
else if (channel ==6'b010001) nextState=ch17;
else if (channel ==6'b010010) nextState=ch18;
else if (channel ==6'b010011) nextState=ch19;
else if (channel ==6'b010100) nextState=ch20;
else if (channel ==6'b010101) nextState=ch21;
else if (channel ==6'b010110) nextState=ch22;
else if (channel ==6'b010111) nextState=ch23;
else if (channel ==6'b011000) nextState=ch24;
else if (channel ==6'b011001) nextState=ch25;
else if (channel ==6'b011010) nextState=ch26;
else if (channel ==6'b011011) nextState=ch27;
else if (channel ==6'b011100) nextState=ch28;
else if (channel ==6'b011101) nextState=ch29;
else if (channel ==6'b011110) nextState=ch30;
else if (channel ==6'b011111) nextState=ch31;
else if (channel ==6'b100000) nextState=ch32;
else if (channel ==6'b100001) nextState=ch33;
else if (channel ==6'b100010) nextState=ch34;
else if (channel ==6'b100011) nextState=ch35;
else if (channel ==6'b100100) nextState=ch36;
else if (channel ==6'b100101) nextState=ch37;
else if (channel ==6'b100110) nextState=ch38;
else if (channel ==6'b100111) nextState=ch39;
else if (channel ==6'b101000) nextState=ch40;
else if (channel ==6'b101001) nextState=ch41;
else if (channel ==6'b101010) nextState=ch42;
else if (channel ==6'b101011) nextState=ch43;
else if (channel ==6'b101100) nextState=ch44;
else if (channel ==6'b101101) nextState=ch45;
else if (channel ==6'b101110) nextState=ch46;
else if (channel ==6'b101111) nextState=ch47;
else if (channel ==6'b110000) nextState=ch48;
else if (channel ==6'b110001) nextState=ch49;
else if (channel ==6'b110010) nextState=ch50;
else if (channel ==6'b110011) nextState=ch51;
else if (channel ==6'b110100) nextState=ch52;
else if (channel ==6'b000000) nextState=ch0;
else if (channel ==6'b110110) nextState=ch54;
else if (channel ==6'b110111) nextState=ch55;
else if (channel ==6'b111000) nextState=ch56;
else if (channel ==6'b111001) nextState=ch57;
else if (channel ==6'b111010) nextState=ch58;
else if (channel ==6'b111011) nextState=ch59;
else if (channel ==6'b111100) nextState=ch60;
else if (channel ==6'b111101) nextState=ch61;
else if (channel ==6'b111110) nextState=ch62;
else nextState=ch63;

ch54: 
if (channel == 6'b110110) nextState=ch54;
else if (channel ==6'b000001) nextState=ch1;
else if (channel ==6'b000010) nextState=ch2;
else if (channel ==6'b000011) nextState=ch3;
else if (channel ==6'b000100) nextState=ch4;
else if (channel ==6'b000101) nextState=ch5;
else if (channel ==6'b000110) nextState=ch6;
else if (channel ==6'b000111) nextState=ch7;
else if (channel ==6'b001000) nextState=ch8;
else if (channel ==6'b001001) nextState=ch9;
else if (channel ==6'b001010) nextState=ch10;
else if (channel ==6'b001011) nextState=ch11;
else if (channel ==6'b001100) nextState=ch12;
else if (channel ==6'b001101) nextState=ch13;
else if (channel ==6'b001110) nextState=ch14;
else if (channel ==6'b001111) nextState=ch15;
else if (channel ==6'b010000) nextState=ch16;
else if (channel ==6'b010001) nextState=ch17;
else if (channel ==6'b010010) nextState=ch18;
else if (channel ==6'b010011) nextState=ch19;
else if (channel ==6'b010100) nextState=ch20;
else if (channel ==6'b010101) nextState=ch21;
else if (channel ==6'b010110) nextState=ch22;
else if (channel ==6'b010111) nextState=ch23;
else if (channel ==6'b011000) nextState=ch24;
else if (channel ==6'b011001) nextState=ch25;
else if (channel ==6'b011010) nextState=ch26;
else if (channel ==6'b011011) nextState=ch27;
else if (channel ==6'b011100) nextState=ch28;
else if (channel ==6'b011101) nextState=ch29;
else if (channel ==6'b011110) nextState=ch30;
else if (channel ==6'b011111) nextState=ch31;
else if (channel ==6'b100000) nextState=ch32;
else if (channel ==6'b100001) nextState=ch33;
else if (channel ==6'b100010) nextState=ch34;
else if (channel ==6'b100011) nextState=ch35;
else if (channel ==6'b100100) nextState=ch36;
else if (channel ==6'b100101) nextState=ch37;
else if (channel ==6'b100110) nextState=ch38;
else if (channel ==6'b100111) nextState=ch39;
else if (channel ==6'b101000) nextState=ch40;
else if (channel ==6'b101001) nextState=ch41;
else if (channel ==6'b101010) nextState=ch42;
else if (channel ==6'b101011) nextState=ch43;
else if (channel ==6'b101100) nextState=ch44;
else if (channel ==6'b101101) nextState=ch45;
else if (channel ==6'b101110) nextState=ch46;
else if (channel ==6'b101111) nextState=ch47;
else if (channel ==6'b110000) nextState=ch48;
else if (channel ==6'b110001) nextState=ch49;
else if (channel ==6'b110010) nextState=ch50;
else if (channel ==6'b110011) nextState=ch51;
else if (channel ==6'b110100) nextState=ch52;
else if (channel ==6'b110101) nextState=ch53;
else if (channel ==6'b000000) nextState=ch0;
else if (channel ==6'b110111) nextState=ch55;
else if (channel ==6'b111000) nextState=ch56;
else if (channel ==6'b111001) nextState=ch57;
else if (channel ==6'b111010) nextState=ch58;
else if (channel ==6'b111011) nextState=ch59;
else if (channel ==6'b111100) nextState=ch60;
else if (channel ==6'b111101) nextState=ch61;
else if (channel ==6'b111110) nextState=ch62;
else nextState=ch63;

ch55: 
if (channel == 6'b110111) nextState=ch55;
else if (channel ==6'b000001) nextState=ch1;
else if (channel ==6'b000010) nextState=ch2;
else if (channel ==6'b000011) nextState=ch3;
else if (channel ==6'b000100) nextState=ch4;
else if (channel ==6'b000101) nextState=ch5;
else if (channel ==6'b000110) nextState=ch6;
else if (channel ==6'b000111) nextState=ch7;
else if (channel ==6'b001000) nextState=ch8;
else if (channel ==6'b001001) nextState=ch9;
else if (channel ==6'b001010) nextState=ch10;
else if (channel ==6'b001011) nextState=ch11;
else if (channel ==6'b001100) nextState=ch12;
else if (channel ==6'b001101) nextState=ch13;
else if (channel ==6'b001110) nextState=ch14;
else if (channel ==6'b001111) nextState=ch15;
else if (channel ==6'b010000) nextState=ch16;
else if (channel ==6'b010001) nextState=ch17;
else if (channel ==6'b010010) nextState=ch18;
else if (channel ==6'b010011) nextState=ch19;
else if (channel ==6'b010100) nextState=ch20;
else if (channel ==6'b010101) nextState=ch21;
else if (channel ==6'b010110) nextState=ch22;
else if (channel ==6'b010111) nextState=ch23;
else if (channel ==6'b011000) nextState=ch24;
else if (channel ==6'b011001) nextState=ch25;
else if (channel ==6'b011010) nextState=ch26;
else if (channel ==6'b011011) nextState=ch27;
else if (channel ==6'b011100) nextState=ch28;
else if (channel ==6'b011101) nextState=ch29;
else if (channel ==6'b011110) nextState=ch30;
else if (channel ==6'b011111) nextState=ch31;
else if (channel ==6'b100000) nextState=ch32;
else if (channel ==6'b100001) nextState=ch33;
else if (channel ==6'b100010) nextState=ch34;
else if (channel ==6'b100011) nextState=ch35;
else if (channel ==6'b100100) nextState=ch36;
else if (channel ==6'b100101) nextState=ch37;
else if (channel ==6'b100110) nextState=ch38;
else if (channel ==6'b100111) nextState=ch39;
else if (channel ==6'b101000) nextState=ch40;
else if (channel ==6'b101001) nextState=ch41;
else if (channel ==6'b101010) nextState=ch42;
else if (channel ==6'b101011) nextState=ch43;
else if (channel ==6'b101100) nextState=ch44;
else if (channel ==6'b101101) nextState=ch45;
else if (channel ==6'b101110) nextState=ch46;
else if (channel ==6'b101111) nextState=ch47;
else if (channel ==6'b110000) nextState=ch48;
else if (channel ==6'b110001) nextState=ch49;
else if (channel ==6'b110010) nextState=ch50;
else if (channel ==6'b110011) nextState=ch51;
else if (channel ==6'b110100) nextState=ch52;
else if (channel ==6'b110101) nextState=ch53;
else if (channel ==6'b110110) nextState=ch54;
else if (channel ==6'b000000) nextState=ch0;
else if (channel ==6'b111000) nextState=ch56;
else if (channel ==6'b111001) nextState=ch57;
else if (channel ==6'b111010) nextState=ch58;
else if (channel ==6'b111011) nextState=ch59;
else if (channel ==6'b111100) nextState=ch60;
else if (channel ==6'b111101) nextState=ch61;
else if (channel ==6'b111110) nextState=ch62;
else nextState=ch63;

ch56: 
if (channel == 6'b111000) nextState=ch56;
else if (channel ==6'b000001) nextState=ch1;
else if (channel ==6'b000010) nextState=ch2;
else if (channel ==6'b000011) nextState=ch3;
else if (channel ==6'b000100) nextState=ch4;
else if (channel ==6'b000101) nextState=ch5;
else if (channel ==6'b000110) nextState=ch6;
else if (channel ==6'b000111) nextState=ch7;
else if (channel ==6'b001000) nextState=ch8;
else if (channel ==6'b001001) nextState=ch9;
else if (channel ==6'b001010) nextState=ch10;
else if (channel ==6'b001011) nextState=ch11;
else if (channel ==6'b001100) nextState=ch12;
else if (channel ==6'b001101) nextState=ch13;
else if (channel ==6'b001110) nextState=ch14;
else if (channel ==6'b001111) nextState=ch15;
else if (channel ==6'b010000) nextState=ch16;
else if (channel ==6'b010001) nextState=ch17;
else if (channel ==6'b010010) nextState=ch18;
else if (channel ==6'b010011) nextState=ch19;
else if (channel ==6'b010100) nextState=ch20;
else if (channel ==6'b010101) nextState=ch21;
else if (channel ==6'b010110) nextState=ch22;
else if (channel ==6'b010111) nextState=ch23;
else if (channel ==6'b011000) nextState=ch24;
else if (channel ==6'b011001) nextState=ch25;
else if (channel ==6'b011010) nextState=ch26;
else if (channel ==6'b011011) nextState=ch27;
else if (channel ==6'b011100) nextState=ch28;
else if (channel ==6'b011101) nextState=ch29;
else if (channel ==6'b011110) nextState=ch30;
else if (channel ==6'b011111) nextState=ch31;
else if (channel ==6'b100000) nextState=ch32;
else if (channel ==6'b100001) nextState=ch33;
else if (channel ==6'b100010) nextState=ch34;
else if (channel ==6'b100011) nextState=ch35;
else if (channel ==6'b100100) nextState=ch36;
else if (channel ==6'b100101) nextState=ch37;
else if (channel ==6'b100110) nextState=ch38;
else if (channel ==6'b100111) nextState=ch39;
else if (channel ==6'b101000) nextState=ch40;
else if (channel ==6'b101001) nextState=ch41;
else if (channel ==6'b101010) nextState=ch42;
else if (channel ==6'b101011) nextState=ch43;
else if (channel ==6'b101100) nextState=ch44;
else if (channel ==6'b101101) nextState=ch45;
else if (channel ==6'b101110) nextState=ch46;
else if (channel ==6'b101111) nextState=ch47;
else if (channel ==6'b110000) nextState=ch48;
else if (channel ==6'b110001) nextState=ch49;
else if (channel ==6'b110010) nextState=ch50;
else if (channel ==6'b110011) nextState=ch51;
else if (channel ==6'b110100) nextState=ch52;
else if (channel ==6'b110101) nextState=ch53;
else if (channel ==6'b110110) nextState=ch54;
else if (channel ==6'b110111) nextState=ch55;
else if (channel ==6'b000000) nextState=ch0;
else if (channel ==6'b111001) nextState=ch57;
else if (channel ==6'b111010) nextState=ch58;
else if (channel ==6'b111011) nextState=ch59;
else if (channel ==6'b111100) nextState=ch60;
else if (channel ==6'b111101) nextState=ch61;
else if (channel ==6'b111110) nextState=ch62;
else nextState=ch63;

ch57: 
if (channel == 6'b111001) nextState=ch57;
else if (channel ==6'b000001) nextState=ch1;
else if (channel ==6'b000010) nextState=ch2;
else if (channel ==6'b000011) nextState=ch3;
else if (channel ==6'b000100) nextState=ch4;
else if (channel ==6'b000101) nextState=ch5;
else if (channel ==6'b000110) nextState=ch6;
else if (channel ==6'b000111) nextState=ch7;
else if (channel ==6'b001000) nextState=ch8;
else if (channel ==6'b001001) nextState=ch9;
else if (channel ==6'b001010) nextState=ch10;
else if (channel ==6'b001011) nextState=ch11;
else if (channel ==6'b001100) nextState=ch12;
else if (channel ==6'b001101) nextState=ch13;
else if (channel ==6'b001110) nextState=ch14;
else if (channel ==6'b001111) nextState=ch15;
else if (channel ==6'b010000) nextState=ch16;
else if (channel ==6'b010001) nextState=ch17;
else if (channel ==6'b010010) nextState=ch18;
else if (channel ==6'b010011) nextState=ch19;
else if (channel ==6'b010100) nextState=ch20;
else if (channel ==6'b010101) nextState=ch21;
else if (channel ==6'b010110) nextState=ch22;
else if (channel ==6'b010111) nextState=ch23;
else if (channel ==6'b011000) nextState=ch24;
else if (channel ==6'b011001) nextState=ch25;
else if (channel ==6'b011010) nextState=ch26;
else if (channel ==6'b011011) nextState=ch27;
else if (channel ==6'b011100) nextState=ch28;
else if (channel ==6'b011101) nextState=ch29;
else if (channel ==6'b011110) nextState=ch30;
else if (channel ==6'b011111) nextState=ch31;
else if (channel ==6'b100000) nextState=ch32;
else if (channel ==6'b100001) nextState=ch33;
else if (channel ==6'b100010) nextState=ch34;
else if (channel ==6'b100011) nextState=ch35;
else if (channel ==6'b100100) nextState=ch36;
else if (channel ==6'b100101) nextState=ch37;
else if (channel ==6'b100110) nextState=ch38;
else if (channel ==6'b100111) nextState=ch39;
else if (channel ==6'b101000) nextState=ch40;
else if (channel ==6'b101001) nextState=ch41;
else if (channel ==6'b101010) nextState=ch42;
else if (channel ==6'b101011) nextState=ch43;
else if (channel ==6'b101100) nextState=ch44;
else if (channel ==6'b101101) nextState=ch45;
else if (channel ==6'b101110) nextState=ch46;
else if (channel ==6'b101111) nextState=ch47;
else if (channel ==6'b110000) nextState=ch48;
else if (channel ==6'b110001) nextState=ch49;
else if (channel ==6'b110010) nextState=ch50;
else if (channel ==6'b110011) nextState=ch51;
else if (channel ==6'b110100) nextState=ch52;
else if (channel ==6'b110101) nextState=ch53;
else if (channel ==6'b110110) nextState=ch54;
else if (channel ==6'b110111) nextState=ch55;
else if (channel ==6'b111000) nextState=ch56;
else if (channel ==6'b000000) nextState=ch0;
else if (channel ==6'b111010) nextState=ch58;
else if (channel ==6'b111011) nextState=ch59;
else if (channel ==6'b111100) nextState=ch60;
else if (channel ==6'b111101) nextState=ch61;
else if (channel ==6'b111110) nextState=ch62;
else nextState=ch63;

ch58: 
if (channel == 6'b111010) nextState=ch58;
else if (channel ==6'b000001) nextState=ch1;
else if (channel ==6'b000010) nextState=ch2;
else if (channel ==6'b000011) nextState=ch3;
else if (channel ==6'b000100) nextState=ch4;
else if (channel ==6'b000101) nextState=ch5;
else if (channel ==6'b000110) nextState=ch6;
else if (channel ==6'b000111) nextState=ch7;
else if (channel ==6'b001000) nextState=ch8;
else if (channel ==6'b001001) nextState=ch9;
else if (channel ==6'b001010) nextState=ch10;
else if (channel ==6'b001011) nextState=ch11;
else if (channel ==6'b001100) nextState=ch12;
else if (channel ==6'b001101) nextState=ch13;
else if (channel ==6'b001110) nextState=ch14;
else if (channel ==6'b001111) nextState=ch15;
else if (channel ==6'b010000) nextState=ch16;
else if (channel ==6'b010001) nextState=ch17;
else if (channel ==6'b010010) nextState=ch18;
else if (channel ==6'b010011) nextState=ch19;
else if (channel ==6'b010100) nextState=ch20;
else if (channel ==6'b010101) nextState=ch21;
else if (channel ==6'b010110) nextState=ch22;
else if (channel ==6'b010111) nextState=ch23;
else if (channel ==6'b011000) nextState=ch24;
else if (channel ==6'b011001) nextState=ch25;
else if (channel ==6'b011010) nextState=ch26;
else if (channel ==6'b011011) nextState=ch27;
else if (channel ==6'b011100) nextState=ch28;
else if (channel ==6'b011101) nextState=ch29;
else if (channel ==6'b011110) nextState=ch30;
else if (channel ==6'b011111) nextState=ch31;
else if (channel ==6'b100000) nextState=ch32;
else if (channel ==6'b100001) nextState=ch33;
else if (channel ==6'b100010) nextState=ch34;
else if (channel ==6'b100011) nextState=ch35;
else if (channel ==6'b100100) nextState=ch36;
else if (channel ==6'b100101) nextState=ch37;
else if (channel ==6'b100110) nextState=ch38;
else if (channel ==6'b100111) nextState=ch39;
else if (channel ==6'b101000) nextState=ch40;
else if (channel ==6'b101001) nextState=ch41;
else if (channel ==6'b101010) nextState=ch42;
else if (channel ==6'b101011) nextState=ch43;
else if (channel ==6'b101100) nextState=ch44;
else if (channel ==6'b101101) nextState=ch45;
else if (channel ==6'b101110) nextState=ch46;
else if (channel ==6'b101111) nextState=ch47;
else if (channel ==6'b110000) nextState=ch48;
else if (channel ==6'b110001) nextState=ch49;
else if (channel ==6'b110010) nextState=ch50;
else if (channel ==6'b110011) nextState=ch51;
else if (channel ==6'b110100) nextState=ch52;
else if (channel ==6'b110101) nextState=ch53;
else if (channel ==6'b110110) nextState=ch54;
else if (channel ==6'b110111) nextState=ch55;
else if (channel ==6'b111000) nextState=ch56;
else if (channel ==6'b111001) nextState=ch57;
else if (channel ==6'b000000) nextState=ch0;
else if (channel ==6'b111011) nextState=ch59;
else if (channel ==6'b111100) nextState=ch60;
else if (channel ==6'b111101) nextState=ch61;
else if (channel ==6'b111110) nextState=ch62;
else nextState=ch63;

ch59: 
if (channel == 6'b111011) nextState=ch59;
else if (channel ==6'b000001) nextState=ch1;
else if (channel ==6'b000010) nextState=ch2;
else if (channel ==6'b000011) nextState=ch3;
else if (channel ==6'b000100) nextState=ch4;
else if (channel ==6'b000101) nextState=ch5;
else if (channel ==6'b000110) nextState=ch6;
else if (channel ==6'b000111) nextState=ch7;
else if (channel ==6'b001000) nextState=ch8;
else if (channel ==6'b001001) nextState=ch9;
else if (channel ==6'b001010) nextState=ch10;
else if (channel ==6'b001011) nextState=ch11;
else if (channel ==6'b001100) nextState=ch12;
else if (channel ==6'b001101) nextState=ch13;
else if (channel ==6'b001110) nextState=ch14;
else if (channel ==6'b001111) nextState=ch15;
else if (channel ==6'b010000) nextState=ch16;
else if (channel ==6'b010001) nextState=ch17;
else if (channel ==6'b010010) nextState=ch18;
else if (channel ==6'b010011) nextState=ch19;
else if (channel ==6'b010100) nextState=ch20;
else if (channel ==6'b010101) nextState=ch21;
else if (channel ==6'b010110) nextState=ch22;
else if (channel ==6'b010111) nextState=ch23;
else if (channel ==6'b011000) nextState=ch24;
else if (channel ==6'b011001) nextState=ch25;
else if (channel ==6'b011010) nextState=ch26;
else if (channel ==6'b011011) nextState=ch27;
else if (channel ==6'b011100) nextState=ch28;
else if (channel ==6'b011101) nextState=ch29;
else if (channel ==6'b011110) nextState=ch30;
else if (channel ==6'b011111) nextState=ch31;
else if (channel ==6'b100000) nextState=ch32;
else if (channel ==6'b100001) nextState=ch33;
else if (channel ==6'b100010) nextState=ch34;
else if (channel ==6'b100011) nextState=ch35;
else if (channel ==6'b100100) nextState=ch36;
else if (channel ==6'b100101) nextState=ch37;
else if (channel ==6'b100110) nextState=ch38;
else if (channel ==6'b100111) nextState=ch39;
else if (channel ==6'b101000) nextState=ch40;
else if (channel ==6'b101001) nextState=ch41;
else if (channel ==6'b101010) nextState=ch42;
else if (channel ==6'b101011) nextState=ch43;
else if (channel ==6'b101100) nextState=ch44;
else if (channel ==6'b101101) nextState=ch45;
else if (channel ==6'b101110) nextState=ch46;
else if (channel ==6'b101111) nextState=ch47;
else if (channel ==6'b110000) nextState=ch48;
else if (channel ==6'b110001) nextState=ch49;
else if (channel ==6'b110010) nextState=ch50;
else if (channel ==6'b110011) nextState=ch51;
else if (channel ==6'b110100) nextState=ch52;
else if (channel ==6'b110101) nextState=ch53;
else if (channel ==6'b110110) nextState=ch54;
else if (channel ==6'b110111) nextState=ch55;
else if (channel ==6'b111000) nextState=ch56;
else if (channel ==6'b111001) nextState=ch57;
else if (channel ==6'b111010) nextState=ch58;
else if (channel ==6'b000000) nextState=ch0;
else if (channel ==6'b111100) nextState=ch60;
else if (channel ==6'b111101) nextState=ch61;
else if (channel ==6'b111110) nextState=ch62;
else nextState=ch63;

ch60: 
if (channel == 6'b111100) nextState=ch60;
else if (channel ==6'b000001) nextState=ch1;
else if (channel ==6'b000010) nextState=ch2;
else if (channel ==6'b000011) nextState=ch3;
else if (channel ==6'b000100) nextState=ch4;
else if (channel ==6'b000101) nextState=ch5;
else if (channel ==6'b000110) nextState=ch6;
else if (channel ==6'b000111) nextState=ch7;
else if (channel ==6'b001000) nextState=ch8;
else if (channel ==6'b001001) nextState=ch9;
else if (channel ==6'b001010) nextState=ch10;
else if (channel ==6'b001011) nextState=ch11;
else if (channel ==6'b001100) nextState=ch12;
else if (channel ==6'b001101) nextState=ch13;
else if (channel ==6'b001110) nextState=ch14;
else if (channel ==6'b001111) nextState=ch15;
else if (channel ==6'b010000) nextState=ch16;
else if (channel ==6'b010001) nextState=ch17;
else if (channel ==6'b010010) nextState=ch18;
else if (channel ==6'b010011) nextState=ch19;
else if (channel ==6'b010100) nextState=ch20;
else if (channel ==6'b010101) nextState=ch21;
else if (channel ==6'b010110) nextState=ch22;
else if (channel ==6'b010111) nextState=ch23;
else if (channel ==6'b011000) nextState=ch24;
else if (channel ==6'b011001) nextState=ch25;
else if (channel ==6'b011010) nextState=ch26;
else if (channel ==6'b011011) nextState=ch27;
else if (channel ==6'b011100) nextState=ch28;
else if (channel ==6'b011101) nextState=ch29;
else if (channel ==6'b011110) nextState=ch30;
else if (channel ==6'b011111) nextState=ch31;
else if (channel ==6'b100000) nextState=ch32;
else if (channel ==6'b100001) nextState=ch33;
else if (channel ==6'b100010) nextState=ch34;
else if (channel ==6'b100011) nextState=ch35;
else if (channel ==6'b100100) nextState=ch36;
else if (channel ==6'b100101) nextState=ch37;
else if (channel ==6'b100110) nextState=ch38;
else if (channel ==6'b100111) nextState=ch39;
else if (channel ==6'b101000) nextState=ch40;
else if (channel ==6'b101001) nextState=ch41;
else if (channel ==6'b101010) nextState=ch42;
else if (channel ==6'b101011) nextState=ch43;
else if (channel ==6'b101100) nextState=ch44;
else if (channel ==6'b101101) nextState=ch45;
else if (channel ==6'b101110) nextState=ch46;
else if (channel ==6'b101111) nextState=ch47;
else if (channel ==6'b110000) nextState=ch48;
else if (channel ==6'b110001) nextState=ch49;
else if (channel ==6'b110010) nextState=ch50;
else if (channel ==6'b110011) nextState=ch51;
else if (channel ==6'b110100) nextState=ch52;
else if (channel ==6'b110101) nextState=ch53;
else if (channel ==6'b110110) nextState=ch54;
else if (channel ==6'b110111) nextState=ch55;
else if (channel ==6'b111000) nextState=ch56;
else if (channel ==6'b111001) nextState=ch57;
else if (channel ==6'b111010) nextState=ch58;
else if (channel ==6'b111011) nextState=ch59;
else if (channel ==6'b111100) nextState=ch60;
else if (channel ==6'b111101) nextState=ch61;
else if (channel ==6'b111110) nextState=ch62;
else nextState=ch63;

ch61: 
if (channel == 6'b111101) nextState=ch61;
else if (channel ==6'b000001) nextState=ch1;
else if (channel ==6'b000010) nextState=ch2;
else if (channel ==6'b000011) nextState=ch3;
else if (channel ==6'b000100) nextState=ch4;
else if (channel ==6'b000101) nextState=ch5;
else if (channel ==6'b000110) nextState=ch6;
else if (channel ==6'b000111) nextState=ch7;
else if (channel ==6'b001000) nextState=ch8;
else if (channel ==6'b001001) nextState=ch9;
else if (channel ==6'b001010) nextState=ch10;
else if (channel ==6'b001011) nextState=ch11;
else if (channel ==6'b001100) nextState=ch12;
else if (channel ==6'b001101) nextState=ch13;
else if (channel ==6'b001110) nextState=ch14;
else if (channel ==6'b001111) nextState=ch15;
else if (channel ==6'b010000) nextState=ch16;
else if (channel ==6'b010001) nextState=ch17;
else if (channel ==6'b010010) nextState=ch18;
else if (channel ==6'b010011) nextState=ch19;
else if (channel ==6'b010100) nextState=ch20;
else if (channel ==6'b010101) nextState=ch21;
else if (channel ==6'b010110) nextState=ch22;
else if (channel ==6'b010111) nextState=ch23;
else if (channel ==6'b011000) nextState=ch24;
else if (channel ==6'b011001) nextState=ch25;
else if (channel ==6'b011010) nextState=ch26;
else if (channel ==6'b011011) nextState=ch27;
else if (channel ==6'b011100) nextState=ch28;
else if (channel ==6'b011101) nextState=ch29;
else if (channel ==6'b011110) nextState=ch30;
else if (channel ==6'b011111) nextState=ch31;
else if (channel ==6'b100000) nextState=ch32;
else if (channel ==6'b100001) nextState=ch33;
else if (channel ==6'b100010) nextState=ch34;
else if (channel ==6'b100011) nextState=ch35;
else if (channel ==6'b100100) nextState=ch36;
else if (channel ==6'b100101) nextState=ch37;
else if (channel ==6'b100110) nextState=ch38;
else if (channel ==6'b100111) nextState=ch39;
else if (channel ==6'b101000) nextState=ch40;
else if (channel ==6'b101001) nextState=ch41;
else if (channel ==6'b101010) nextState=ch42;
else if (channel ==6'b101011) nextState=ch43;
else if (channel ==6'b101100) nextState=ch44;
else if (channel ==6'b101101) nextState=ch45;
else if (channel ==6'b101110) nextState=ch46;
else if (channel ==6'b101111) nextState=ch47;
else if (channel ==6'b110000) nextState=ch48;
else if (channel ==6'b110001) nextState=ch49;
else if (channel ==6'b110010) nextState=ch50;
else if (channel ==6'b110011) nextState=ch51;
else if (channel ==6'b110100) nextState=ch52;
else if (channel ==6'b110101) nextState=ch53;
else if (channel ==6'b110110) nextState=ch54;
else if (channel ==6'b110111) nextState=ch55;
else if (channel ==6'b111000) nextState=ch56;
else if (channel ==6'b111001) nextState=ch57;
else if (channel ==6'b111010) nextState=ch58;
else if (channel ==6'b111011) nextState=ch59;
else if (channel ==6'b111100) nextState=ch60;
else if (channel ==6'b000000) nextState=ch0;
else if (channel ==6'b111110) nextState=ch62;
else nextState=ch63;

ch62: 
if (channel == 6'b111110) nextState=ch62;
else if (channel ==6'b000001) nextState=ch1;
else if (channel ==6'b000010) nextState=ch2;
else if (channel ==6'b000011) nextState=ch3;
else if (channel ==6'b000100) nextState=ch4;
else if (channel ==6'b000101) nextState=ch5;
else if (channel ==6'b000110) nextState=ch6;
else if (channel ==6'b000111) nextState=ch7;
else if (channel ==6'b001000) nextState=ch8;
else if (channel ==6'b001001) nextState=ch9;
else if (channel ==6'b001010) nextState=ch10;
else if (channel ==6'b001011) nextState=ch11;
else if (channel ==6'b001100) nextState=ch12;
else if (channel ==6'b001101) nextState=ch13;
else if (channel ==6'b001110) nextState=ch14;
else if (channel ==6'b001111) nextState=ch15;
else if (channel ==6'b010000) nextState=ch16;
else if (channel ==6'b010001) nextState=ch17;
else if (channel ==6'b010010) nextState=ch18;
else if (channel ==6'b010011) nextState=ch19;
else if (channel ==6'b010100) nextState=ch20;
else if (channel ==6'b010101) nextState=ch21;
else if (channel ==6'b010110) nextState=ch22;
else if (channel ==6'b010111) nextState=ch23;
else if (channel ==6'b011000) nextState=ch24;
else if (channel ==6'b011001) nextState=ch25;
else if (channel ==6'b011010) nextState=ch26;
else if (channel ==6'b011011) nextState=ch27;
else if (channel ==6'b011100) nextState=ch28;
else if (channel ==6'b011101) nextState=ch29;
else if (channel ==6'b011110) nextState=ch30;
else if (channel ==6'b011111) nextState=ch31;
else if (channel ==6'b100000) nextState=ch32;
else if (channel ==6'b100001) nextState=ch33;
else if (channel ==6'b100010) nextState=ch34;
else if (channel ==6'b100011) nextState=ch35;
else if (channel ==6'b100100) nextState=ch36;
else if (channel ==6'b100101) nextState=ch37;
else if (channel ==6'b100110) nextState=ch38;
else if (channel ==6'b100111) nextState=ch39;
else if (channel ==6'b101000) nextState=ch40;
else if (channel ==6'b101001) nextState=ch41;
else if (channel ==6'b101010) nextState=ch42;
else if (channel ==6'b101011) nextState=ch43;
else if (channel ==6'b101100) nextState=ch44;
else if (channel ==6'b101101) nextState=ch45;
else if (channel ==6'b101110) nextState=ch46;
else if (channel ==6'b101111) nextState=ch47;
else if (channel ==6'b110000) nextState=ch48;
else if (channel ==6'b110001) nextState=ch49;
else if (channel ==6'b110010) nextState=ch50;
else if (channel ==6'b110011) nextState=ch51;
else if (channel ==6'b110100) nextState=ch52;
else if (channel ==6'b110101) nextState=ch53;
else if (channel ==6'b110110) nextState=ch54;
else if (channel ==6'b110111) nextState=ch55;
else if (channel ==6'b111000) nextState=ch56;
else if (channel ==6'b111001) nextState=ch57;
else if (channel ==6'b111010) nextState=ch58;
else if (channel ==6'b111011) nextState=ch59;
else if (channel ==6'b111100) nextState=ch60;
else if (channel ==6'b111101) nextState=ch61;
else if (channel ==6'b000000) nextState=ch0;
else nextState=ch63;


ch63:if (channel ==6'b111111) nextState=ch63;
else nextState = ch0;

default: nextState = ch0;
endcase
assign channel_op = channel;
//(currentState==ch0 | currentState==ch1 |currentState==ch2 | currentState==ch3 |currentState==ch4 | currentState==ch5 | currentState==ch6 | currentState==ch7 | currentState==ch8 | currentState==ch9 | currentState==ch10 | currentState==ch11 | currentState==ch12 | currentState==ch13 | currentState==ch14 | currentState==ch15 | currentState==ch16 | currentState==ch17 | currentState==ch18 | currentState==ch19 | currentState==ch20 | currentState==ch21 | currentState==ch22 | currentState==ch23 | currentState==ch24 | currentState==ch25 | currentState==ch26 | currentState==ch27 | currentState==ch28 | currentState==ch29 | currentState==ch30 | currentState==ch31);
assign data_op = data;
assign concat_data1=reg1+reg2;

// Read and write fifo pointers (We put -2, because on the case of DEPTH=8
    // clog2(DEPTH) = 3, then 1:0, 2 bits, we count from 0 to 3
     reg [(clogb2(DEPTH)-1):0] rd_ptr, wr_ptr;
	  
	  
    // Declare the fifo memory (RAM that allow read and write at the same time)
    // reg [7:0] [3:0], create an array of 4 elements of 8 bits
    reg [(NUM_BITS-1):0] fifo_mem[(DEPTH-1):0];
    
    
    // Combinational part that calculate the empty/full flags
    assign empty = (fifo_counter==0);
    assign full = (fifo_counter==DEPTH);

    
    // Sequential circuit that will handle the fifo_counter, which is used to 
    // detect if the fifo is empty or full.
    always @(posedge clk or negedge rst_n)
    begin

        if (~rst_n)
            fifo_counter = 0;
        else if( (!full && wr_en1) && ( !empty && rd_en1 ) ) 
            fifo_counter = fifo_counter;     // If read and write don't change counter          
        else if (!full && wr_en1)  
            fifo_counter = fifo_counter + 1; // Only write increment            
        else if (!empty && rd_en1)  
            fifo_counter = fifo_counter - 1; // Only read decrement                                          
    end
    
    // Sequential circuit to handle reading on the fifo
    always @( posedge clk or negedge rst_n)
    begin
        if( ~rst_n )
            fifo_out = 0;
        else
            begin
              // Give some data if not empty and we want to read
              if ( !empty && rd_en1 )
                begin
                    fifo_out = fifo_mem[rd_ptr];
                    // synthesis translate_off                    
                    $display("Popping value: %d at %t",fifo_mem[rd_ptr],$time);                    
                    // synthesis translate_on
                end                    
                                 
                                                       
            end
    end
    
    // Sequential circuit to handle writing to the fifo
    always @(posedge clk)
    begin    
       if (!full && wr_en1)
        begin
            fifo_mem[ wr_ptr ] = fifo_in;
            // synthesis translate_off                    
            $display("Pushing value: %d at %t",fifo_in,$time);                    
            // synthesis translate_on
        end                            
    end
    
    // Sequential circut to handle the read/write pointers
    always@(posedge clk or negedge rst_n)
    begin
        if( ~rst_n )
        begin
            // In the beginning the pointers are the same
            wr_ptr = 0;
            rd_ptr = 0;
        end
        else
        begin
            // We're not full and someone want to write, so we increment the write pointer
            if( !full && wr_en1 )
                wr_ptr = wr_ptr + 1;              
            
            // We're not empty and someone want to read, so we decrement the read pointer
            if( !empty && rd_en1 )
                rd_ptr = rd_ptr + 1;          
        end    
    end    	 
	 
	 function integer clogb2;
    input [31:0] depth;
        begin
            depth = depth - 1;
            for(clogb2=0; depth>0; clogb2=clogb2+1)
                depth = depth >> 1;
        end
    endfunction
	 
endmodule


